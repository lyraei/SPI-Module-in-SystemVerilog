select_slave = 2;
send_request = 1;
             // AAAAAAAA0BBBBBBBB0PPPP000000 
send_data = 28'b1111111101100110000001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011000100110000011000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0001100101011000100100000000;
expected_data = 28'b1111101110100000000000000000;
@(next_data);

send_data = 28'b1110001100101010100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0011011100110010000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010001101101101000111000000;
expected_data = 28'b0110111010000000000000000000;
@(next_data);

send_data = 28'b1010010000111000001000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b0101000001111110101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001001001010101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011101011101100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011111000101010000001000000;
expected_data = 28'b1100001010100000000000000000;
@(next_data);

send_data = 28'b1111001001100111100010000000;
expected_data = 28'b0111111000000000000000000000;
@(next_data);

send_data = 28'b1110011000100011000011000000;
expected_data = 28'b0111100110000000000000000000;
@(next_data);

send_data = 28'b0111010100101000000100000000;
expected_data = 28'b1011100110100000000000000000;
@(next_data);

send_data = 28'b0001010001001101100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0111101100001101100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101000011100100111000000;
expected_data = 28'b1111011000100000000000000000;
@(next_data);

send_data = 28'b1010100101001011001000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1010110001010100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000011000100101001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011010000111111000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100101000100111000001000000;
expected_data = 28'b1011001000100000000000000000;
@(next_data);

send_data = 28'b1100011100000010100010000000;
expected_data = 28'b0100111000000000000000000000;
@(next_data);

send_data = 28'b0001111000000000000011000000;
expected_data = 28'b0110001100000000000000000000;
@(next_data);

send_data = 28'b0010011100101000000100000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0011101000101110000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0001001101101101000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111010000100011100111000000;
expected_data = 28'b0010011010000000000000000000;
@(next_data);

send_data = 28'b1001000001011001001000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b1010001100100100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110001100111110001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100001100001000000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111101100010010000001000000;
expected_data = 28'b0101001100000000000000000000;
@(next_data);

send_data = 28'b0011111000111110100010000000;
expected_data = 28'b0111111110000000000000000000;
@(next_data);

send_data = 28'b0010010100010100000011000000;
expected_data = 28'b0001111110000000000000000000;
@(next_data);

send_data = 28'b1001000000100001100100000000;
expected_data = 28'b1101111110100000000000000000;
@(next_data);

send_data = 28'b1100011000100011000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1001000100000011100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011111100001111000111000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b1101000001111001101000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0010111001101101001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101000100001000101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001011100001100100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001010001010110100001000000;
expected_data = 28'b0011000000000000000000000000;
@(next_data);

send_data = 28'b1000110000101011000010000000;
expected_data = 28'b1011110100100000000000000000;
@(next_data);

send_data = 28'b1000110001010010000011000000;
expected_data = 28'b0100011010000000000000000000;
@(next_data);

send_data = 28'b1110100001010111100100000000;
expected_data = 28'b0111101100000000000000000000;
@(next_data);

send_data = 28'b1100011001011111000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1110001001000000000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110001000001010000111000000;
expected_data = 28'b1100010010100000000000000000;
@(next_data);

send_data = 28'b1011011000111111001000000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1101111000000111101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001000110010101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110100000011110100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111010100111101000001000000;
expected_data = 28'b1010010100100000000000000000;
@(next_data);

send_data = 28'b0011110100010101000010000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1111110001001001000011000000;
expected_data = 28'b0001111000000000000000000000;
@(next_data);

send_data = 28'b0011111000001010000100000000;
expected_data = 28'b0110111100000000000000000000;
@(next_data);