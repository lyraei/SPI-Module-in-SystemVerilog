select_slave = 0;
send_request = 1;

send_data = 28'b0000000000000000000000000000;
expected_data = '0;
@(next_data);

send_data = 28'b0000000000011100000001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000011000101110000010000000;
expected_data = 28'b0011100000000000000000000000;
@(next_data);

send_data = 28'b1100111001100011100011000000;
expected_data = 28'b1111101100010000000000000000;
@(next_data);

send_data = 28'b1100011001111001100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100001100101111100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100011101000100100110000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0111111000100010100111000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0101110101001000101000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0110111001000111101001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b0011110001100100101010000000;
expected_data = 28'b0110111000000000000000000000;
@(next_data);

send_data = 28'b1110001101101110001011000000;
expected_data = 28'b0011110001000000000000000000;
@(next_data);

send_data = 28'b0010110000101111101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0001000101101000101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000000001101000101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111111100011000101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110011000100101000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001010100010010100001000000;
expected_data = 28'b0001110000000000000000000000;
@(next_data);

send_data = 28'b0001011101010100100010000000;
expected_data = 28'b1011000000010000000000000000;
@(next_data);

send_data = 28'b1100001101001011100011000000;
expected_data = 28'b1111111000010000000000000000;
@(next_data);

send_data = 28'b1001110001111011000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000000000010100000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010011100110111000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000010101010100000111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b1010010001110111001000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001100101001110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1001100001110101101010000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b1100101101011100001011000000;
expected_data = 28'b1110100001010000000000000000;
@(next_data);

send_data = 28'b1110010101011000101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0110011101100111001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000101100010000001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011100010111001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000000101010001100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001100001110000000001000000;
expected_data = 28'b0101111000000000000000000000;
@(next_data);

send_data = 28'b0011011101001011100010000000;
expected_data = 28'b0111100001000000000000000000;
@(next_data);

send_data = 28'b1010010101011111100011000000;
expected_data = 28'b1110100001010000000000000000;
@(next_data);

send_data = 28'b1110001001101100100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100010001110101000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010001001010110100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111111100111110000111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010001001100101101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000110100000100001001000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b1011111101010101101010000000;
expected_data = 28'b0000110100000000000000000000;
@(next_data);

send_data = 28'b1011000001101001001011000000;
expected_data = 28'b1100000100010000000000000000;
@(next_data);

send_data = 28'b1101101001110010001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0010001000011110001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110011101100011001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100100000101110001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101101110110000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010011100011100000001000000;
expected_data = 28'b1101111100010000000000000000;
@(next_data);

send_data = 28'b1011001101111111000010000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b0101110001001101100011000000;
expected_data = 28'b0100110101000000000000000000;
@(next_data);

send_data = 28'b1110011000101101100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111001100000001000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011101001110000000110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0111110101000110100111000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0011110001000100001000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001100111111001001000000;
expected_data = 28'b0000101001000000000000000000;
@(next_data);

send_data = 28'b1010100100001111001010000000;
expected_data = 28'b1100110100010000000000000000;
@(next_data);

send_data = 28'b1000100000010011001011000000;
expected_data = 28'b1101011101010000000000000000;
@(next_data);

send_data = 28'b0100011101011010001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1111001001101010001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100000100001011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101101010001101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001010100000000000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111011001011010100001000000;
expected_data = 28'b1001010101010000000000000000;
@(next_data);

send_data = 28'b1010111100011000000010000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b1110011101100001100011000000;
expected_data = 28'b1101111100010000000000000000;
@(next_data);

send_data = 28'b1101000000011011000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011001000010100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100100100001001100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1010001001110000100111000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0011000000111100001000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0000111000110001001001000000;
expected_data = 28'b0000101001000000000000000000;
@(next_data);

send_data = 28'b1010011101101000101010000000;
expected_data = 28'b0000111000000000000000000000;
@(next_data);

send_data = 28'b0101110101110011001011000000;
expected_data = 28'b1101100100010000000000000000;
@(next_data);

send_data = 28'b0011111101101010101100000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0001111000000011001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010001001101111101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111001100010001001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000100101011000100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101001101001011000001000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b1010100101111010100010000000;
expected_data = 28'b1100010101010000000000000000;
@(next_data);

send_data = 28'b0101111100000011000011000000;
expected_data = 28'b0101111000000000000000000000;
@(next_data);

send_data = 28'b1010000100001100000100000000;
expected_data = 28'b1100000001010000000000000000;
@(next_data);

send_data = 28'b0001001100100001000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000001001100111100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1010111101011001100111000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0001010001110110001000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011011001100111001001000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b0110001001100100001010000000;
expected_data = 28'b1100101001010000000000000000;
@(next_data);

send_data = 28'b0101010000111110001011000000;
expected_data = 28'b0110001000000000000000000000;
@(next_data);

send_data = 28'b1010111101111001101100000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1000011001111111001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110011100101111001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101000011010001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010100001100100000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010001001101001100001000000;
expected_data = 28'b1110000000010000000000000000;
@(next_data);

send_data = 28'b0111010101000111000010000000;
expected_data = 28'b1111000100010000000000000000;
@(next_data);

send_data = 28'b1111010000110100000011000000;
expected_data = 28'b1111101100010000000000000000;
@(next_data);

send_data = 28'b0011000001010101000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100001101011110000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111000100001000100110000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b1111100000111100000111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101011000010011101000000000;
expected_data = 28'b0000001101000000000000000000;
@(next_data);

send_data = 28'b1101110001001011101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1101101001000000101010000000;
expected_data = 28'b1010010000010000000000000000;
@(next_data);

send_data = 28'b1010100101000101101011000000;
expected_data = 28'b1010011001010000000000000000;
@(next_data);

send_data = 28'b0101100001011000101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1010000001001101101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100011100101001001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111000100110100001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100110100000100000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110001000001101100001000000;
expected_data = 28'b1100010101010000000000000000;
@(next_data);

send_data = 28'b0100000001011010000010000000;
expected_data = 28'b1111100101010000000000000000;
@(next_data);

send_data = 28'b1110111100010101000011000000;
expected_data = 28'b1111111101110000000000000000;
@(next_data);

send_data = 28'b0010110001000110000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101000011001100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111011100101001000110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1110110101101110100111000000;
expected_data = 28'b0000001101000000000000000000;
@(next_data);

send_data = 28'b0011101000110100101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100101000100100101001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b0110100001111000101010000000;
expected_data = 28'b0100101000000000000000000000;
@(next_data);

send_data = 28'b1011000101110111001011000000;
expected_data = 28'b0110100000000000000000000000;
@(next_data);

send_data = 28'b1101100101010110001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0111101100111100001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101001001110110001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011010001000011001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010100100010101000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010011001101011000001000000;
expected_data = 28'b0111111100000000000000000000;
@(next_data);

send_data = 28'b1000111001001100000010000000;
expected_data = 28'b0111000000000000000000000000;
@(next_data);

send_data = 28'b1010111101100001000011000000;
expected_data = 28'b0111011101000000000000000000;
@(next_data);

send_data = 28'b0001110100101010100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011010001001101000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100111101000000000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001001001100010100111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110000001110100001000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0110000100010010101001000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b1011110101000010001010000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b1101100001011011001011000000;
expected_data = 28'b1100001101010000000000000000;
@(next_data);

send_data = 28'b1010001100111100001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1011111101110011001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110110101101011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011010001001000001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100010101110000000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001110100010001100001000000;
expected_data = 28'b0110010101000000000000000000;
@(next_data);

send_data = 28'b0011110001110001100010000000;
expected_data = 28'b0011111000000000000000000000;
@(next_data);

send_data = 28'b1010110101101110100011000000;
expected_data = 28'b1101111100010000000000000000;
@(next_data);

send_data = 28'b0110001101001011000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100001101010000100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000110100000001000110000000;
expected_data = 28'b0000001101000000000000000000;
@(next_data);

send_data = 28'b0000100000100111000111000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0011110001101000101000000000;
expected_data = 28'b0000001101000000000000000000;
@(next_data);

send_data = 28'b0001100100010100001001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1110001000001111101010000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b1010000100010111001011000000;
expected_data = 28'b1001111000010000000000000000;
@(next_data);

send_data = 28'b0000001101010000001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1010110001110111001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101011100011011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001110001011110101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000010001101010100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000101101101100100001000000;
expected_data = 28'b1010111101010000000000000000;
@(next_data);

send_data = 28'b0111111001011011100010000000;
expected_data = 28'b0101001000000000000000000000;
@(next_data);

send_data = 28'b0111100000110001100011000000;
expected_data = 28'b1100100101010000000000000000;
@(next_data);

send_data = 28'b0011010101101011000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001001001010101100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001101001011011100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1000001001100101100111000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1001110000100101001000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0000010100000010101001000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b0011011000010000001010000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1010100101101100101011000000;
expected_data = 28'b0011011001000000000000000000;
@(next_data);

send_data = 28'b0001110001010100001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0001011100101001001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010100001010011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010110100111111001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001111101010101000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100111101000100000001000000;
expected_data = 28'b0111010100000000000000000000;
@(next_data);

send_data = 28'b1110001101010101000010000000;
expected_data = 28'b0100011101000000000000000000;
@(next_data);

send_data = 28'b1011101000111000100011000000;
expected_data = 28'b0101110100000000000000000000;
@(next_data);

send_data = 28'b1010010001001011000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100010101101011100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011100101111010100110000000;
expected_data = 28'b0000001101000000000000000000;
@(next_data);

send_data = 28'b0101000101100101000111000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0010011000111000101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100110100010100001001000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b0111010000101101101010000000;
expected_data = 28'b0100110101000000000000000000;
@(next_data);

send_data = 28'b1010010000111000101011000000;
expected_data = 28'b0111010001000000000000000000;
@(next_data);

send_data = 28'b1110101000000110101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0111000101000101101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100110100011100001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100001100111101101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010100001111100100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101110000111100000001000000;
expected_data = 28'b1010111101010000000000000000;
@(next_data);

send_data = 28'b0100110101101000000010000000;
expected_data = 28'b0010010001000000000000000000;
@(next_data);

send_data = 28'b0011001000101111100011000000;
expected_data = 28'b1011111100010000000000000000;
@(next_data);

send_data = 28'b1001011100100110100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001011101111101000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011001000110100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0101101000000111000111000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1101100000101110001000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b1011001001011010001001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1010101000001111001010000000;
expected_data = 28'b1100111000010000000000000000;
@(next_data);

send_data = 28'b0101111101110100001011000000;
expected_data = 28'b1101011000010000000000000000;
@(next_data);

send_data = 28'b0100000100100001001100000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1100000001100101101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000110100111011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100111101001010101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000100000101010000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100000001010011100001000000;
expected_data = 28'b0011010000000000000000000000;
@(next_data);

send_data = 28'b1111101101011000100010000000;
expected_data = 28'b1110011101010000000000000000;
@(next_data);

send_data = 28'b1011100001011101000011000000;
expected_data = 28'b0100111001000000000000000000;
@(next_data);

send_data = 28'b1100110100110101100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101110001010000100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111001001100010000110000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b1001101101001010000111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b1000011100001100101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000111001000010101001000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b0100001100010110101010000000;
expected_data = 28'b1111001000010000000000000000;
@(next_data);

send_data = 28'b1011110100110100101011000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b1100110101011010001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1010010001111101101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000100000110011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101001110010001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000000100100010100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010000001100111000001000000;
expected_data = 28'b1011110000010000000000000000;
@(next_data);

send_data = 28'b0111111100100110100010000000;
expected_data = 28'b1110111001010000000000000000;
@(next_data);

send_data = 28'b0011110100100101000011000000;
expected_data = 28'b1011001001010000000000000000;
@(next_data);

send_data = 28'b1101111100101100100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111110100001001000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100100100101101000110000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0010101001001000100111000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110000101010111101000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b1101001000010110101001000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1111111101100010101010000000;
expected_data = 28'b1010111000010000000000000000;
@(next_data);

send_data = 28'b1011101000101011001011000000;
expected_data = 28'b1000000101010000000000000000;
@(next_data);

send_data = 28'b0001000001100011001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0101010001011110001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011001101000000101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000100101011100101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010110100100111000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011101000101101100001000000;
expected_data = 28'b1101111100010000000000000000;
@(next_data);

send_data = 28'b1100100000001111000010000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b1100100000000110000011000000;
expected_data = 28'b1111011100010000000000000000;
@(next_data);

send_data = 28'b0011101100111011000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111111100100101000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010110101000010100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0011011000111000000111000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0110101100001101001000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0000011101111100101001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1111011001001101101010000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0110110000100101101011000000;
expected_data = 28'b1000101000010000000000000000;
@(next_data);

send_data = 28'b0110100001101001101100000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1001111100110100101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101111001011100101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001010001001110001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111111001110100100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110001000111011000001000000;
expected_data = 28'b0001010100000000000000000000;
@(next_data);

send_data = 28'b0001101000001010000010000000;
expected_data = 28'b0001010001000000000000000000;
@(next_data);

send_data = 28'b0111101100011011100011000000;
expected_data = 28'b1110111100010000000000000000;
@(next_data);

send_data = 28'b0010101100001100100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111110100000000000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001100001111010100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000010101101011100111000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1000010000101000101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100111001110110001001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1001101001101110001010000000;
expected_data = 28'b0100111001000000000000000000;
@(next_data);

send_data = 28'b1111111000001100001011000000;
expected_data = 28'b1110011000010000000000000000;
@(next_data);

send_data = 28'b0000011100011000101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110110000001001001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010111100111101101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100111000100111001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011110101000011100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011101111111100001000000;
expected_data = 28'b1011011000010000000000000000;
@(next_data);

send_data = 28'b0001001001001100100010000000;
expected_data = 28'b1111100000010000000000000000;
@(next_data);

send_data = 28'b1000110100011100100011000000;
expected_data = 28'b1110111100010000000000000000;
@(next_data);

send_data = 28'b1100110001001010000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010101001001111100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101111101101000100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1111010101010000100111000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0110000100100000101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110000101100000101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1011001100010110101010000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b1011010001100100101011000000;
expected_data = 28'b1100110100010000000000000000;
@(next_data);

send_data = 28'b1111100100010101101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011101101000000101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010010101010100001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010000101100011001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000101101001010000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010110001000110100001000000;
expected_data = 28'b1111011100010000000000000000;
@(next_data);

send_data = 28'b1010010001000110100010000000;
expected_data = 28'b1010000100010000000000000000;
@(next_data);

send_data = 28'b0100111001011100100011000000;
expected_data = 28'b0111101101000000000000000000;
@(next_data);

send_data = 28'b0001100000010111000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101000000100111000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010101001011011100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111110001110010000111000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b0001000001101001001000000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b1001000001110101101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0110000101010101001010000000;
expected_data = 28'b1111000001010000000000000000;
@(next_data);

send_data = 28'b1110101001010000001011000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b0010001000000010101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0010001100011011101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001011101001110001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000111100011011001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110001100111000000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111000000110111100001000000;
expected_data = 28'b1111001101010000000000000000;
@(next_data);

send_data = 28'b0001110000100101000010000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b0010011101001011000011000000;
expected_data = 28'b1111011100010000000000000000;
@(next_data);

send_data = 28'b1101110100010011100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101010001110101000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111110101011111000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010100001110101100111000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b0111011001110000001000000000;
expected_data = 28'b0000001101000000000000000000;
@(next_data);

send_data = 28'b1100010101001011101001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b0001110101110101001010000000;
expected_data = 28'b1011101101010000000000000000;
@(next_data);

send_data = 28'b0001010100001100001011000000;
expected_data = 28'b0001110101000000000000000000;
@(next_data);

send_data = 28'b0011111001111101101100000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b1101001000110111001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011001100010101001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001100000011001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001011100111010100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011101010110100001000000;
expected_data = 28'b1010001000010000000000000000;
@(next_data);

send_data = 28'b0010000101010000000010000000;
expected_data = 28'b1010101001010000000000000000;
@(next_data);

send_data = 28'b1001011101110010100011000000;
expected_data = 28'b1101111100010000000000000000;
@(next_data);

send_data = 28'b1100010001011011100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011000100000100000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001100111010100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010000000011110000111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101000100100001001000000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1000001001010100001001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1011100101111100101010000000;
expected_data = 28'b1111111000010000000000000000;
@(next_data);

send_data = 28'b1100000101110001001011000000;
expected_data = 28'b1100011100010000000000000000;
@(next_data);

send_data = 28'b1110000000100000101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0001000000001011101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111111101001110101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011111001101011001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100111101111011100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011111000000011100001000000;
expected_data = 28'b1101100001010000000000000000;
@(next_data);

send_data = 28'b1010110101101100000010000000;
expected_data = 28'b1011100100010000000000000000;
@(next_data);

send_data = 28'b0011100001111011000011000000;
expected_data = 28'b0111011101000000000000000000;
@(next_data);

send_data = 28'b0100110000000110100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111100101111011000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111111001110010000110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1010000101001001000111000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0011011101100010101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101111001011100001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0101110000101101101010000000;
expected_data = 28'b1010001000010000000000000000;
@(next_data);

send_data = 28'b1001001001110101001011000000;
expected_data = 28'b0101110001000000000000000000;
@(next_data);

send_data = 28'b0111001100000001001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011110101101110001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101101011011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111101100111111101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000111000011110100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111110001111001100001000000;
expected_data = 28'b0101000100000000000000000000;
@(next_data);

send_data = 28'b0001011101011010000010000000;
expected_data = 28'b0000111101000000000000000000;
@(next_data);

send_data = 28'b1011100000100110100011000000;
expected_data = 28'b1110101101010000000000000000;
@(next_data);

send_data = 28'b1100110100101001100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101100001011101000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110100101000100100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000001001110001000111000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b1001011000011000001000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b1000110000001110001001000000;
expected_data = 28'b0000101001000000000000000000;
@(next_data);

send_data = 28'b1000011100000111001010000000;
expected_data = 28'b1111010000010000000000000000;
@(next_data);

send_data = 28'b0100010000101001001011000000;
expected_data = 28'b1111100101010000000000000000;
@(next_data);

send_data = 28'b0011110100110001101100000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0100111100001111001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111111001011010001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100110100001000101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010111001000110000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011110001010000100001000000;
expected_data = 28'b1010001000010000000000000000;
@(next_data);

send_data = 28'b0000101000110101100010000000;
expected_data = 28'b0001110101000000000000000000;
@(next_data);

send_data = 28'b1110000101010110000011000000;
expected_data = 28'b1111010101010000000000000000;
@(next_data);

send_data = 28'b0111011001010011100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001000100001000000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101011100101101100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001000101100000111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b1011001000100000001000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b1101010001101111101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0001010001000011001010000000;
expected_data = 28'b1010110001010000000000000000;
@(next_data);

send_data = 28'b1010110000111010001011000000;
expected_data = 28'b0001010001000000000000000000;
@(next_data);

send_data = 28'b0101100001000000001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1101011001111011001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111010100100011101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010110001101010101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101111100001101100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001010001111100100001000000;
expected_data = 28'b0100010001000000000000000000;
@(next_data);

send_data = 28'b1000110001011000000010000000;
expected_data = 28'b0110110100000000000000000000;
@(next_data);

send_data = 28'b1001001000000011000011000000;
expected_data = 28'b0111111100000000000000000000;
@(next_data);

send_data = 28'b0100111100010000100100000000;
expected_data = 28'b1000000010010000000000000000;
@(next_data);

send_data = 28'b0111111100110111100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000001001100100100110000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1011011000101100100111000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1010101101010101101000000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b1001100001100010001001000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0011001001011000101010000000;
expected_data = 28'b1110100001010000000000000000;
@(next_data);

send_data = 28'b1011010101110001001011000000;
expected_data = 28'b0011001000000000000000000000;
@(next_data);

send_data = 28'b1011100000110110001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1111100000011011001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010100101001101001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010110000100101101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010110000001111000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001001001101000001000000;
expected_data = 28'b1000111001010000000000000000;
@(next_data);

send_data = 28'b1111100101010101000010000000;
expected_data = 28'b0010100001000000000000000000;
@(next_data);

send_data = 28'b1100010001000101100011000000;
expected_data = 28'b0101011100000000000000000000;
@(next_data);

send_data = 28'b0011100101101001000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001010100000001100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111110101011101000110000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0010110001000001000111000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0111010100010000001000000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0101000100100011001001000000;
expected_data = 28'b0000101001000000000000000000;
@(next_data);

send_data = 28'b0110101101111001101010000000;
expected_data = 28'b0101000100000000000000000000;
@(next_data);

send_data = 28'b0110010000110100001011000000;
expected_data = 28'b0110101100000000000000000000;
@(next_data);

send_data = 28'b0010100000011010001100000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0111010100110100001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101011000101000101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111011000010101101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111011001011111000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101001101110000001000000;
expected_data = 28'b1011100001010000000000000000;
@(next_data);

send_data = 28'b0000011001111110000010000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1000011101010001000011000000;
expected_data = 28'b1111101100010000000000000000;
@(next_data);

send_data = 28'b1110100101100001000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101111101011001000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011001001000110100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0100101101010011000111000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b1101111000100010001000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001000001001101001001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1001111100010101001010000000;
expected_data = 28'b0001000010000000000000000000;
@(next_data);

send_data = 28'b1101010100000011101011000000;
expected_data = 28'b1110000101010000000000000000;
@(next_data);

send_data = 28'b0100110101101101101100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1010010101100110001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001010101000011001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100110100110011001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111100000001110100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110101001100110100001000000;
expected_data = 28'b1101101101010000000000000000;
@(next_data);

send_data = 28'b1011111101011110100010000000;
expected_data = 28'b1010011100010000000000000000;
@(next_data);

send_data = 28'b0000001101110100100011000000;
expected_data = 28'b0100001001000000000000000000;
@(next_data);

send_data = 28'b1111000101111000000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000000000001101000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110010100001100100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110000101101001000111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b1000110001011010101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111111001010101101001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b0000011001010101001010000000;
expected_data = 28'b0111111001000000000000000000;
@(next_data);

send_data = 28'b0011110001111101101011000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1010001000101111001100000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b0111011000101110101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101001101100110001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000101100010010101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100001000101011000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101011100011011000001000000;
expected_data = 28'b1110110000010000000000000000;
@(next_data);

send_data = 28'b1000100100111111100010000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b0111100000011010100011000000;
expected_data = 28'b1111011001010000000000000000;
@(next_data);

send_data = 28'b1011100000101010000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011001101001000000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011000101010110000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101001100100101100111000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1111110100000100101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101110100001110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011001000100000101010000000;
expected_data = 28'b1010001101010000000000000000;
@(next_data);

send_data = 28'b1110010101011010001011000000;
expected_data = 28'b0011001000000000000000000000;
@(next_data);

send_data = 28'b0111101101011000001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0110111101100101101101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101100000010111101110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010001001100011101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011111000111100100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010111001001011000001000000;
expected_data = 28'b1100010101010000000000000000;
@(next_data);

send_data = 28'b0010000100100101100010000000;
expected_data = 28'b1011100001010000000000000000;
@(next_data);

send_data = 28'b0011111101001011100011000000;
expected_data = 28'b1111111000010000000000000000;
@(next_data);

send_data = 28'b0111111001101111100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101100010000100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000011000000111100110000000;
expected_data = 28'b0000001101000000000000000000;
@(next_data);

send_data = 28'b0010000101000110100111000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b1000011001100111101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000010100100100001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0000110000011001001010000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b0011010101101111101011000000;
expected_data = 28'b0000110001000000000000000000;
@(next_data);

send_data = 28'b0000001101011110101100000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1011000001000000001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100000100011000001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001110001110011001111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010111101001001000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001010100010001100001000000;
expected_data = 28'b0001110101000000000000000000;
@(next_data);

send_data = 28'b1001110001010001000010000000;
expected_data = 28'b0011011001000000000000000000;
@(next_data);

send_data = 28'b1100011100101001100011000000;
expected_data = 28'b0111111100000000000000000000;
@(next_data);

send_data = 28'b0101101000111100000100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001101001001100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001000111111100110000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1110000100100110000111000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0101010101000101101000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110100100100001101001000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1101001100011110001010000000;
expected_data = 28'b0110100101000000000000000000;
@(next_data);

send_data = 28'b1010011100101110101011000000;
expected_data = 28'b1010110100010000000000000000;
@(next_data);

send_data = 28'b0011111000110101001100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1111000001001111001101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000011101100110001110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001110000101000101111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010111001010000100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100011101100111100001000000;
expected_data = 28'b1000110101010000000000000000;
@(next_data);

send_data = 28'b0110011000111110000010000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1001100101110100100011000000;
expected_data = 28'b1001101100010000000000000000;
@(next_data);

send_data = 28'b0011101101111111100100000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110111100000000000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110001101101010100000000000;
expected_data = 28'b0110111101000000000000000000;
@(next_data);

send_data = 28'b1011001101100000000000000000;
expected_data = 28'b1000111001010000000000000000;
@(next_data);

send_data = 28'b0111011000110111100000000000;
expected_data = 28'b1111001101010000000000000000;
@(next_data);

send_data = 28'b1011110000001000000001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1101100100010000100001000000;
expected_data = 28'b1010110001010000000000000000;
@(next_data);

send_data = 28'b1001001101101000100001000000;
expected_data = 28'b1111100000010000000000000000;
@(next_data);

send_data = 28'b0100100100000100100001000000;
expected_data = 28'b0100001001000000000000000000;
@(next_data);

send_data = 28'b1001000100111111100010000000;
expected_data = 28'b0100000010000000000000000000;
@(next_data);

send_data = 28'b1111111001111011100010000000;
expected_data = 28'b1110111001010000000000000000;
@(next_data);

send_data = 28'b0111010101101110000010000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b0001000100010110000010000000;
expected_data = 28'b1010101100010000000000000000;
@(next_data);

send_data = 28'b1010001001001110000011000000;
expected_data = 28'b1111111101110000000000000000;
@(next_data);

send_data = 28'b0011111100000000100011000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100010000000001000011000000;
expected_data = 28'b0111111001000000000000000000;
@(next_data);

send_data = 28'b0100101100000001100011000000;
expected_data = 28'b0001000010000000000000000000;
@(next_data);

send_data = 28'b0101010100000000000100000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b0000111100000000100100000000;
expected_data = 28'b0101010101000000000000000000;
@(next_data);

send_data = 28'b1110101100000001000100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0100110000000001100100000000;
expected_data = 28'b0011101001000000000000000000;
@(next_data);

send_data = 28'b0001100100000000000101000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b1100011100110101100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101101000010000101000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0010110101011001100101000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b0000000101001110100111000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0001000001110011000111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001000000101110100111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b0010000000001010100111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b0000100000100001001000000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b0011001000011100001000000000;
expected_data = 28'b0000110100000000000000000000;
@(next_data);

send_data = 28'b0001011001010111001000000000;
expected_data = 28'b0000101001000000000000000000;
@(next_data);

send_data = 28'b0110011101111001101000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1000010100111111101001000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1101010000101001001001000000;
expected_data = 28'b1111101100010000000000000000;
@(next_data);

send_data = 28'b1111011101011001101001000000;
expected_data = 28'b1010110001010000000000000000;
@(next_data);

send_data = 28'b1011010000000100001001000000;
expected_data = 28'b1000100100010000000000000000;
@(next_data);

send_data = 28'b0010111100110011001010000000;
expected_data = 28'b1100110001010000000000000000;
@(next_data);

send_data = 28'b1010110100100011101010000000;
expected_data = 28'b0010111100000000000000000000;
@(next_data);

send_data = 28'b1001111000000110101010000000;
expected_data = 28'b1101001100010000000000000000;
@(next_data);

send_data = 28'b1101000001101011001010000000;
expected_data = 28'b1110001001010000000000000000;
@(next_data);

send_data = 28'b0100110100100100001011000000;
expected_data = 28'b1011000000010000000000000000;
@(next_data);

send_data = 28'b1001100100110101001011000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0101010000001000101011000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110101101111000001011000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1001101001011101001011000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1000001001100100100101000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1000001000010100100110000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0001001000111101100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001001000110101100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1100101101010010100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101100111010100110000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011010101111011000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);