select_slave = 1;
send_request = 1;

send_data = 28'b0000000000000000000000000000;
expected_data = 28'b0010111100000000000000000000;
@(next_data);

send_data = 28'b0000000000011100000001000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011000101110000010000000;
expected_data = 28'b0011100000000000000000000000;
@(next_data);

send_data = 28'b1100111001100011100011000000;
expected_data = 28'b0010010100000000000000000000;
@(next_data);

send_data = 28'b1100011001111001100100000000;
expected_data = 28'b0110011100000000000000000000;
@(next_data);

send_data = 28'b1100001100101111100101000000;
expected_data = 28'b1000110001000000000000000000;
@(next_data);

send_data = 28'b0100011101000100100110000000;
expected_data = 28'b1010001001000000000000000000;
@(next_data);

send_data = 28'b0111111000100010100111000000;
expected_data = 28'b0100011100000000000000000000;
@(next_data);

send_data = 28'b0101110101001000101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0110111001000111101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0011110001100100101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110001101101110001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010110000101111101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000101101000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000001101000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111100011000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110011000100101000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001010100010010100001000000;
expected_data = 28'b1011000001000000000000000000;
@(next_data);

send_data = 28'b0001011101010100100010000000;
expected_data = 28'b1011000001000000000000000000;
@(next_data);

send_data = 28'b1100001101001011100011000000;
expected_data = 28'b0100000100000000000000000000;
@(next_data);

send_data = 28'b1001110001111011000100000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b0000000000010100000101000000;
expected_data = 28'b0011100000000000000000000000;
@(next_data);

send_data = 28'b1010011100110111000110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000010101010100000111000000;
expected_data = 28'b1101100101000000000000000000;
@(next_data);

send_data = 28'b1010010001110111001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001100101001110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1001100001110101101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1100101101011100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110010101011000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110011101100111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000101100010000001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011100010111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000101010001100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001100001110000000001000000;
expected_data = 28'b1010010001000000000000000000;
@(next_data);

send_data = 28'b0011011101001011100010000000;
expected_data = 28'b0111100000000000000000000000;
@(next_data);

send_data = 28'b1010010101011111100011000000;
expected_data = 28'b0101111100000000000000000000;
@(next_data);

send_data = 28'b1110001001101100100100000000;
expected_data = 28'b0101001000000000000000000000;
@(next_data);

send_data = 28'b0100010001110101000101000000;
expected_data = 28'b1100010001000000000000000000;
@(next_data);

send_data = 28'b1010001001010110100110000000;
expected_data = 28'b0110011000000000000000000000;
@(next_data);

send_data = 28'b1111111100111110000111000000;
expected_data = 28'b1101111001000000000000000000;
@(next_data);

send_data = 28'b0010001001100101101000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0000110100000100001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1011111101010101101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011000001101001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101101001110010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010001000011110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110011101100011001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100100000101110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100101101110110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010011100011100000001000000;
expected_data = 28'b1011011101010000000000000000;
@(next_data);

send_data = 28'b1011001101111111000010000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b0101110001001101100011000000;
expected_data = 28'b1011001001000000000000000000;
@(next_data);

send_data = 28'b1110011000101101100100000000;
expected_data = 28'b0010111000000000000000000000;
@(next_data);

send_data = 28'b0111001100000001000101000000;
expected_data = 28'b1100110001000000000000000000;
@(next_data);

send_data = 28'b1011101001110000000110000000;
expected_data = 28'b0100101000000000000000000000;
@(next_data);

send_data = 28'b0111110101000110100111000000;
expected_data = 28'b1100011001000000000000000000;
@(next_data);

send_data = 28'b0011110001000100001000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b1011001100111111001001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1010100100001111001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1000100000010011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0100011101011010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111001001101010001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100000100001011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101101010001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001010100000000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011001011010100001000000;
expected_data = 28'b1001010101000000000000000000;
@(next_data);

send_data = 28'b1010111100011000000010000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b1110011101100001100011000000;
expected_data = 28'b0110000000000000000000000000;
@(next_data);

send_data = 28'b1101000000011011000100000000;
expected_data = 28'b0111001100000000000000000000;
@(next_data);

send_data = 28'b0000011001000010100101000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b1100100100001001100110000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1010001001110000100111000000;
expected_data = 28'b1011011101000000000000000000;
@(next_data);

send_data = 28'b0011000000111100001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0000111000110001001001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1010011101101000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0101110101110011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0011111101101010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111000000011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010001001101111101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111001100010001001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000100101011000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101001101001011000001000000;
expected_data = 28'b1011101001000000000000000000;
@(next_data);

send_data = 28'b1010100101111010100010000000;
expected_data = 28'b1100010101000000000000000000;
@(next_data);

send_data = 28'b0101111100000011000011000000;
expected_data = 28'b1010001101000000000000000000;
@(next_data);

send_data = 28'b1010000100001100000100000000;
expected_data = 28'b0010111100000000000000000000;
@(next_data);

send_data = 28'b0001001100100001000101000000;
expected_data = 28'b0100001000000000000000000000;
@(next_data);

send_data = 28'b0000001001100111100110000000;
expected_data = 28'b0001101000000000000000000000;
@(next_data);

send_data = 28'b1010111101011001100111000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0001010001110110001000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b1011011001100111001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0110001001100100001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0101010000111110001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1010111101111001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011001111111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110011100101111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101000011010001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100001100100000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010001001101001100001000000;
expected_data = 28'b0111000000010000000000000000;
@(next_data);

send_data = 28'b0111010101000111000010000000;
expected_data = 28'b1111000101000000000000000000;
@(next_data);

send_data = 28'b1111010000110100000011000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0011000001010101000100000000;
expected_data = 28'b0111101000000000000000000000;
@(next_data);

send_data = 28'b0100001101011110000101000000;
expected_data = 28'b0110000000000000000000000000;
@(next_data);

send_data = 28'b1111000100001000100110000000;
expected_data = 28'b0110001000000000000000000000;
@(next_data);

send_data = 28'b1111100000111100000111000000;
expected_data = 28'b1000111101000000000000000000;
@(next_data);

send_data = 28'b1101011000010011101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101110001001011101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1101101001000000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010100101000101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101100001011000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010000001001101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100011100101001001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111000100110100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100110100000100000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110001000001101100001000000;
expected_data = 28'b1101010101000000000000000000;
@(next_data);

send_data = 28'b0100000001011010000010000000;
expected_data = 28'b1111100101000000000000000000;
@(next_data);

send_data = 28'b1110111100010101000011000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0010110001000110000100000000;
expected_data = 28'b0111011100000000000000000000;
@(next_data);

send_data = 28'b1101101000011001100101000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b0111011100101001000110000000;
expected_data = 28'b1011011101000000000000000000;
@(next_data);

send_data = 28'b1110110101101110100111000000;
expected_data = 28'b0111011100000000000000000000;
@(next_data);

send_data = 28'b0011101000110100101000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b0100101000100100101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0110100001111000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011000101110111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101100101010110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111101100111100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101001001110110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011010001000011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100100010101000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010011001101011000001000000;
expected_data = 28'b1101001101000000000000000000;
@(next_data);

send_data = 28'b1000111001001100000010000000;
expected_data = 28'b0111000000000000000000000000;
@(next_data);

send_data = 28'b1010111101100001000011000000;
expected_data = 28'b1110100101000000000000000000;
@(next_data);

send_data = 28'b0001110100101010100100000000;
expected_data = 28'b0101011100000000000000000000;
@(next_data);

send_data = 28'b1011010001001101000101000000;
expected_data = 28'b0011101000000000000000000000;
@(next_data);

send_data = 28'b1100111101000000000110000000;
expected_data = 28'b1110111001000000000000000000;
@(next_data);

send_data = 28'b0001001001100010100111000000;
expected_data = 28'b1011000101000000000000000000;
@(next_data);

send_data = 28'b1110000001110100001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0110000100010010101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1011110101000010001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101100001011011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1010001100111100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011111101110011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110110101101011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011010001001000001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100010101110000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001110100010001100001000000;
expected_data = 28'b0010010100010000000000000000;
@(next_data);

send_data = 28'b0011110001110001100010000000;
expected_data = 28'b0011111000000000000000000000;
@(next_data);

send_data = 28'b1010110101101110100011000000;
expected_data = 28'b0010000000100000000000000000;
@(next_data);

send_data = 28'b0110001101001011000100000000;
expected_data = 28'b0101011000000000000000000000;
@(next_data);

send_data = 28'b0100001101010000100101000000;
expected_data = 28'b1100011001000000000000000000;
@(next_data);

send_data = 28'b1000110100000001000110000000;
expected_data = 28'b0110001000000000000000000000;
@(next_data);

send_data = 28'b0000100000100111000111000000;
expected_data = 28'b1111001101000000000000000000;
@(next_data);

send_data = 28'b0011110001101000101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001100100010100001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1110001000001111101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010000100010111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000001101010000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110001110111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101011100011011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001110001011110101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000010001101010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000101101101100100001000000;
expected_data = 28'b0101100100010000000000000000;
@(next_data);

send_data = 28'b0111111001011011100010000000;
expected_data = 28'b0101001000000000000000000000;
@(next_data);

send_data = 28'b0111100000110001100011000000;
expected_data = 28'b0011011000000000000000000000;
@(next_data);

send_data = 28'b0011010101101011000100000000;
expected_data = 28'b0011110000000000000000000000;
@(next_data);

send_data = 28'b1001001001010101100101000000;
expected_data = 28'b0110101000000000000000000000;
@(next_data);

send_data = 28'b1001101001011011100110000000;
expected_data = 28'b1101101101000000000000000000;
@(next_data);

send_data = 28'b1000001001100101100111000000;
expected_data = 28'b1110011001000000000000000000;
@(next_data);

send_data = 28'b1001110000100101001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0000010100000010101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0011011000010000001010000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b1010100101101100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0001110001010100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011100101001001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010100001010011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110100111111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111101010101000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100111101000100000001000000;
expected_data = 28'b1100100101000000000000000000;
@(next_data);

send_data = 28'b1110001101010101000010000000;
expected_data = 28'b0100011100000000000000000000;
@(next_data);

send_data = 28'b1011101000111000100011000000;
expected_data = 28'b1011011001000000000000000000;
@(next_data);

send_data = 28'b1010010001001011000100000000;
expected_data = 28'b0101110100000000000000000000;
@(next_data);

send_data = 28'b0100010101101011100101000000;
expected_data = 28'b0100100000000000000000000000;
@(next_data);

send_data = 28'b0011100101111010100110000000;
expected_data = 28'b0110011100000000000000000000;
@(next_data);

send_data = 28'b0101000101100101000111000000;
expected_data = 28'b0011100100000000000000000000;
@(next_data);

send_data = 28'b0010011000111000101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0100110100010100001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0111010000101101101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010010000111000101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110101000000110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111000101000101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100110100011100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100001100111101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100001111100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101110000111100000001000000;
expected_data = 28'b1010000101010000000000000000;
@(next_data);

send_data = 28'b0100110101101000000010000000;
expected_data = 28'b0010010000000000000000000000;
@(next_data);

send_data = 28'b0011001000101111100011000000;
expected_data = 28'b0110001000000000000000000000;
@(next_data);

send_data = 28'b1001011100100110100100000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b1001011101111101000101000000;
expected_data = 28'b0010111000000000000000000000;
@(next_data);

send_data = 28'b0000011001000110100110000000;
expected_data = 28'b1101110001000000000000000000;
@(next_data);

send_data = 28'b0101101000000111000111000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1101100000101110001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1011001001011010001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1010101000001111001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0101111101110100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0100000100100001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100000001100101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110100111011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100111101001010101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100000101010000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100000001010011100001000000;
expected_data = 28'b1101110001000000000000000000;
@(next_data);

send_data = 28'b1111101101011000100010000000;
expected_data = 28'b1110011101000000000000000000;
@(next_data);

send_data = 28'b1011100001011101000011000000;
expected_data = 28'b1011010101000000000000000000;
@(next_data);

send_data = 28'b1100110100110101100100000000;
expected_data = 28'b0101110000000000000000000000;
@(next_data);

send_data = 28'b0101110001010000100101000000;
expected_data = 28'b1001101001000000000000000000;
@(next_data);

send_data = 28'b1111001001100010000110000000;
expected_data = 28'b0111001000000000000000000000;
@(next_data);

send_data = 28'b1001101101001010000111000000;
expected_data = 28'b1000111001000000000000000000;
@(next_data);

send_data = 28'b1000011100001100101000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1000111001000010101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0100001100010110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011110100110100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1100110101011010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010001111101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000100000110011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101001110010001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000100100010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010000001100111000001000000;
expected_data = 28'b0100011000000000000000000000;
@(next_data);

send_data = 28'b0111111100100110100010000000;
expected_data = 28'b1110111001000000000000000000;
@(next_data);

send_data = 28'b0011110100100101000011000000;
expected_data = 28'b1100110101000000000000000000;
@(next_data);

send_data = 28'b1101111100101100100100000000;
expected_data = 28'b0001111000000000000000000000;
@(next_data);

send_data = 28'b1111110100001001000101000000;
expected_data = 28'b1011111001000000000000000000;
@(next_data);

send_data = 28'b0100100100101101000110000000;
expected_data = 28'b1000001101000000000000000000;
@(next_data);

send_data = 28'b0010101001001000100111000000;
expected_data = 28'b0100100100000000000000000000;
@(next_data);

send_data = 28'b1110000101010111101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1101001000010110101001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1111111101100010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011101000101011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0001000001100011001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101010001011110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011001101000000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000100101011100101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110100100111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101000101101100001000000;
expected_data = 28'b0111101100000000000000000000;
@(next_data);

send_data = 28'b1100100000001111000010000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b1100100000000110000011000000;
expected_data = 28'b0010100100000000000000000000;
@(next_data);

send_data = 28'b0011101100111011000100000000;
expected_data = 28'b0110010000000000000000000000;
@(next_data);

send_data = 28'b0111111100100101000101000000;
expected_data = 28'b0111011000000000000000000000;
@(next_data);

send_data = 28'b1010110101000010100110000000;
expected_data = 28'b0100000000100000000000000000;
@(next_data);

send_data = 28'b0011011000111000000111000000;
expected_data = 28'b1101001101000000000000000000;
@(next_data);

send_data = 28'b0110101100001101001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011101111100101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1111011001001101101010000000;
expected_data = 28'b0111111100000000000000000000;
@(next_data);

send_data = 28'b0110110000100101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0110100001101001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001111100110100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101111001011100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010001001110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111001110100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110001000111011000001000000;
expected_data = 28'b1110011101010000000000000000;
@(next_data);

send_data = 28'b0001101000001010000010000000;
expected_data = 28'b0001010000000000000000000000;
@(next_data);

send_data = 28'b0111101100011011100011000000;
expected_data = 28'b1111000101000000000000000000;
@(next_data);

send_data = 28'b0010101100001100100100000000;
expected_data = 28'b0011110100000000000000000000;
@(next_data);

send_data = 28'b0111110100000000000101000000;
expected_data = 28'b0101011000000000000000000000;
@(next_data);

send_data = 28'b0001100001111010100110000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b0000010101101011100111000000;
expected_data = 28'b0001100000000000000000000000;
@(next_data);

send_data = 28'b1000010000101000101000000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b0100111001110110001001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1001101001101110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1111111000001100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000011100011000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110110000001001001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010111100111101101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100111000100111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011110101000011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011101111111100001000000;
expected_data = 28'b1100010001000000000000000000;
@(next_data);

send_data = 28'b0001001001001100100010000000;
expected_data = 28'b1111100001000000000000000000;
@(next_data);

send_data = 28'b1000110100011100100011000000;
expected_data = 28'b0111010000000000000000000000;
@(next_data);

send_data = 28'b1100110001001010000100000000;
expected_data = 28'b0100011000000000000000000000;
@(next_data);

send_data = 28'b0010101001001111100101000000;
expected_data = 28'b1001100001000000000000000000;
@(next_data);

send_data = 28'b1101111101101000100110000000;
expected_data = 28'b0011111100000000000000000000;
@(next_data);

send_data = 28'b1111010101010000100111000000;
expected_data = 28'b1010000101000000000000000000;
@(next_data);

send_data = 28'b0110000100100000101000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0110000101100000101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1011001100010110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011010001100100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111100100010101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101101000000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010101010100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010000101100011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000101101001010000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110001000110100001000000;
expected_data = 28'b0001111100010000000000000000;
@(next_data);

send_data = 28'b1010010001000110100010000000;
expected_data = 28'b1010000101000000000000000000;
@(next_data);

send_data = 28'b0100111001011100100011000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b0001100000010111000100000000;
expected_data = 28'b0010011100000000000000000000;
@(next_data);

send_data = 28'b0101000000100111000101000000;
expected_data = 28'b0011000000000000000000000000;
@(next_data);

send_data = 28'b1010101001011011100110000000;
expected_data = 28'b0111100000000000000000000000;
@(next_data);

send_data = 28'b0111110001110010000111000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b0001000001101001001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001000001110101101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0110000101010101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110101001010000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010001000000010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010001100011011101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011101001110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000111100011011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110001100111000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111000000110111100001000000;
expected_data = 28'b1101001101000000000000000000;
@(next_data);

send_data = 28'b0001110000100101000010000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b0010011101001011000011000000;
expected_data = 28'b1010100101000000000000000000;
@(next_data);

send_data = 28'b1101110100010011100100000000;
expected_data = 28'b0001001100000000000000000000;
@(next_data);

send_data = 28'b0101010001110101000101000000;
expected_data = 28'b1011101001000000000000000000;
@(next_data);

send_data = 28'b0111110101011111000110000000;
expected_data = 28'b0111111000000000000000000000;
@(next_data);

send_data = 28'b0010100001110101100111000000;
expected_data = 28'b0111110100000000000000000000;
@(next_data);

send_data = 28'b0111011001110000001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100010101001011101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0001110101110101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0001010100001100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0011111001111101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101001000110111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011001100010101001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011001100000011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011100111010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011101010110100001000000;
expected_data = 28'b1000110001000000000000000000;
@(next_data);

send_data = 28'b0010000101010000000010000000;
expected_data = 28'b1010101001000000000000000000;
@(next_data);

send_data = 28'b1001011101110010100011000000;
expected_data = 28'b0111111000000000000000000000;
@(next_data);

send_data = 28'b1100010001011011100100000000;
expected_data = 28'b0100101100000000000000000000;
@(next_data);

send_data = 28'b0011000100000100000101000000;
expected_data = 28'b1000100001000000000000000000;
@(next_data);

send_data = 28'b1011001100111010100110000000;
expected_data = 28'b0010100100000000000000000000;
@(next_data);

send_data = 28'b1010000000011110000111000000;
expected_data = 28'b1100110101000000000000000000;
@(next_data);

send_data = 28'b0101000100100001001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000001001010100001001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1011100101111100101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1100000101110001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110000000100000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000000001011101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111101001110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011111001101011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100111101111011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011111000000011100001000000;
expected_data = 28'b1100011001010000000000000000;
@(next_data);

send_data = 28'b1010110101101100000010000000;
expected_data = 28'b1011100101000000000000000000;
@(next_data);

send_data = 28'b0011100001111011000011000000;
expected_data = 28'b1000101001000000000000000000;
@(next_data);

send_data = 28'b0100110000000110100100000000;
expected_data = 28'b0001110000000000000000000000;
@(next_data);

send_data = 28'b0111100101111011000101000000;
expected_data = 28'b1001100001000000000000000000;
@(next_data);

send_data = 28'b1111111001110010000110000000;
expected_data = 28'b0100010100000000000000000000;
@(next_data);

send_data = 28'b1010000101001001000111000000;
expected_data = 28'b1000001001000000000000000000;
@(next_data);

send_data = 28'b0011011101100010101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1101111001011100001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0101110000101101101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1001001001110101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111001100000001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011110101101110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101101011011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111101100111111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000111000011110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111110001111001100001000000;
expected_data = 28'b1100101101000000000000000000;
@(next_data);

send_data = 28'b0001011101011010000010000000;
expected_data = 28'b0000111100000000000000000000;
@(next_data);

send_data = 28'b1011100000100110100011000000;
expected_data = 28'b0101110000000000000000000000;
@(next_data);

send_data = 28'b1100110100101001100100000000;
expected_data = 28'b0101110000000000000000000000;
@(next_data);

send_data = 28'b0101100001011101000101000000;
expected_data = 28'b1001101001000000000000000000;
@(next_data);

send_data = 28'b0110100101000100100110000000;
expected_data = 28'b0111010000000000000000000000;
@(next_data);

send_data = 28'b0000001001110001000111000000;
expected_data = 28'b0110100100000000000000000000;
@(next_data);

send_data = 28'b1001011000011000001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1000110000001110001001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1000011100000111001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0100010000101001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0011110100110001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111100001111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111111001011010001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100110100001000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010111001000110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011110001010000100001000000;
expected_data = 28'b1011101001000000000000000000;
@(next_data);

send_data = 28'b0000101000110101100010000000;
expected_data = 28'b0001110100000000000000000000;
@(next_data);

send_data = 28'b1110000101010110000011000000;
expected_data = 28'b1001111001000000000000000000;
@(next_data);

send_data = 28'b0111011001010011100100000000;
expected_data = 28'b0111000000000000000000000000;
@(next_data);

send_data = 28'b1001000100001000000101000000;
expected_data = 28'b1110110001000000000000000000;
@(next_data);

send_data = 28'b0101011100101101100110000000;
expected_data = 28'b1101100101000000000000000000;
@(next_data);

send_data = 28'b1011001000101100000111000000;
expected_data = 28'b0101011100000000000000000000;
@(next_data);

send_data = 28'b1011001000100000001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101010001101111101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0001010001000011001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010110000111010001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101100001000000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101011001111011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111010100100011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110001101010101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101111100001101100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001010001111100100001000000;
expected_data = 28'b0111101000000000000000000000;
@(next_data);

send_data = 28'b1000110001011000000010000000;
expected_data = 28'b0110110100000000000000000000;
@(next_data);

send_data = 28'b1001001000000011000011000000;
expected_data = 28'b1100001101000000000000000000;
@(next_data);

send_data = 28'b0100111100010000100100000000;
expected_data = 28'b0100100100000000000000000000;
@(next_data);

send_data = 28'b0111111100110111100101000000;
expected_data = 28'b1001111001000000000000000000;
@(next_data);

send_data = 28'b1000001001100100100110000000;
expected_data = 28'b0100000000100000000000000000;
@(next_data);

send_data = 28'b1011011000101100100111000000;
expected_data = 28'b1111111001000000000000000000;
@(next_data);

send_data = 28'b1010101101010101101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1001100001100010001001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0011001001011000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011010101110001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1011100000110110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111100000011011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100101001101001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110000100101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110000001111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011001001001101000001000000;
expected_data = 28'b1100101001000000000000000000;
@(next_data);

send_data = 28'b1111100101010101000010000000;
expected_data = 28'b0010100000000000000000000000;
@(next_data);

send_data = 28'b1100010001000101100011000000;
expected_data = 28'b1010110001000000000000000000;
@(next_data);

send_data = 28'b0011100101101001000100000000;
expected_data = 28'b0110001000000000000000000000;
@(next_data);

send_data = 28'b0001010100000001100101000000;
expected_data = 28'b0111001000000000000000000000;
@(next_data);

send_data = 28'b1111110101011101000110000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b0010110001000001000111000000;
expected_data = 28'b1000001101000000000000000000;
@(next_data);

send_data = 28'b0111010100010000001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101000100100011001001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b0110101101111001101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0110010000110100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010100000011010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111010100110100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101011000101000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011000010101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111011001011111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101001101110000001000000;
expected_data = 28'b0011010000010000000000000000;
@(next_data);

send_data = 28'b0000011001111110000010000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1000011101010001000011000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1110100101100001000100000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b1101111101011001000101000000;
expected_data = 28'b1101001001000000000000000000;
@(next_data);

send_data = 28'b0011001001000110100110000000;
expected_data = 28'b1011000001000000000000000000;
@(next_data);

send_data = 28'b0100101101010011000111000000;
expected_data = 28'b0011001000000000000000000000;
@(next_data);

send_data = 28'b1101111000100010001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0001000001001101001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1001111100010101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101010100000011101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0100110101101101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010101100110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010101000011001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100110100110011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111100000001110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110101001100110100001000000;
expected_data = 28'b0001010100010000000000000000;
@(next_data);

send_data = 28'b1011111101011110100010000000;
expected_data = 28'b1010011101000000000000000000;
@(next_data);

send_data = 28'b0000001101110100100011000000;
expected_data = 28'b1111110101000000000000000000;
@(next_data);

send_data = 28'b1111000101111000000100000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b0000000000001101000101000000;
expected_data = 28'b1110001001000000000000000000;
@(next_data);

send_data = 28'b1110010100001100100110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110000101101001000111000000;
expected_data = 28'b1001101101000000000000000000;
@(next_data);

send_data = 28'b1000110001011010101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0111111001010101101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0000011001010101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0011110001111101101011000000;
expected_data = 28'b0010000000100000000000000000;
@(next_data);

send_data = 28'b1010001000101111001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111011000101110101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101001101100110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000101100010010101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100001000101011000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101011100011011000001000000;
expected_data = 28'b1001100001000000000000000000;
@(next_data);

send_data = 28'b1000100100111111100010000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b0111100000011010100011000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1011100000101010000100000000;
expected_data = 28'b0011110000000000000000000000;
@(next_data);

send_data = 28'b0011001101001000000101000000;
expected_data = 28'b0111000000000000000000000000;
@(next_data);

send_data = 28'b0011000101010110000110000000;
expected_data = 28'b0010101000000000000000000000;
@(next_data);

send_data = 28'b1101001100100101100111000000;
expected_data = 28'b0011000100000000000000000000;
@(next_data);

send_data = 28'b1111110100000100101000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1101110100001110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011001000100000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110010101011010001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111101101011000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110111101100101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100000010111101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010001001100011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011111000111100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010111001001011000001000000;
expected_data = 28'b1011011101000000000000000000;
@(next_data);

send_data = 28'b0010000100100101100010000000;
expected_data = 28'b1011100001000000000000000000;
@(next_data);

send_data = 28'b0011111101001011100011000000;
expected_data = 28'b1001010101000000000000000000;
@(next_data);

send_data = 28'b0111111001101111100100000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b1100101100010000100101000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b1000011000000111100110000000;
expected_data = 28'b1010111001000000000000000000;
@(next_data);

send_data = 28'b0010000101000110100111000000;
expected_data = 28'b1111101001000000000000000000;
@(next_data);

send_data = 28'b1000011001100111101000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0000010100100100001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0000110000011001001010000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b0011010101101111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000001101011110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011000001000000001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100000100011000001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001110001110011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010111101001001000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010100010001100001000000;
expected_data = 28'b0100000100010000000000000000;
@(next_data);

send_data = 28'b1001110001010001000010000000;
expected_data = 28'b0011011000000000000000000000;
@(next_data);

send_data = 28'b1100011100101001100011000000;
expected_data = 28'b1100000101000000000000000000;
@(next_data);

send_data = 28'b0101101000111100000100000000;
expected_data = 28'b0110001100000000000000000000;
@(next_data);

send_data = 28'b1011001101001001100101000000;
expected_data = 28'b1011010001000000000000000000;
@(next_data);

send_data = 28'b1011001000111111100110000000;
expected_data = 28'b1110101001000000000000000000;
@(next_data);

send_data = 28'b1110000100100110000111000000;
expected_data = 28'b1100111001000000000000000000;
@(next_data);

send_data = 28'b0101010101000101101000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0110100100100001101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1101001100011110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010011100101110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0011111000110101001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111000001001111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011101100110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001110000101000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010111001010000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100011101100111100001000000;
expected_data = 28'b1100111101000000000000000000;
@(next_data);

send_data = 28'b0110011000111110000010000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1001100101110100100011000000;
expected_data = 28'b1110010101000000000000000000;
@(next_data);

send_data = 28'b0011101101111111100100000000;
expected_data = 28'b0100110000000000000000000000;
@(next_data);

send_data = 28'b0110111100110001100101000000;
expected_data = 28'b0111011000000000000000000000;
@(next_data);

send_data = 28'b1101010101011001100110000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b1100000000111011000111000000;
expected_data = 28'b1010101101000000000000000000;
@(next_data);

send_data = 28'b0110111101011110001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000001101100101001000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0010000101001001101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101000100100100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000100101001000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111111101111111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011100111010101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101110000001000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110001010001000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001110000011111100001000000;
expected_data = 28'b1100111001000000000000000000;
@(next_data);

send_data = 28'b0100010000100101100010000000;
expected_data = 28'b1010001101000000000000000000;
@(next_data);

send_data = 28'b0101010100000111100011000000;
expected_data = 28'b1111000001000000000000000000;
@(next_data);

send_data = 28'b1110101100100110000100000000;
expected_data = 28'b0010101000000000000000000000;
@(next_data);

send_data = 28'b0001100101100011100101000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b0110101101101101100110000000;
expected_data = 28'b0001010100000000000000000000;
@(next_data);

send_data = 28'b1000010000010110100111000000;
expected_data = 28'b0110101100000000000000000000;
@(next_data);

send_data = 28'b1011001101101100001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1001110101000110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110011001110010001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0101110101111010101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0001010100000100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100001000011001001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011100000001011001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010111000110011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111001101000010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111111101101010000001000000;
expected_data = 28'b0111100000010000000000000000;
@(next_data);

send_data = 28'b0101001001111011100010000000;
expected_data = 28'b1010101101000000000000000000;
@(next_data);

send_data = 28'b1011001101011010000011000000;
expected_data = 28'b0101101000000000000000000000;
@(next_data);

send_data = 28'b0000100000010111100100000000;
expected_data = 28'b0101100100000000000000000000;
@(next_data);

send_data = 28'b0110011001010110100101000000;
expected_data = 28'b0001000000100000000000000000;
@(next_data);

send_data = 28'b0100011101001111000110000000;
expected_data = 28'b0101010100000000000000000000;
@(next_data);

send_data = 28'b0000110101101000000111000000;
expected_data = 28'b0100011100000000000000000000;
@(next_data);

send_data = 28'b1101011000100110101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100100001001100101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0110101000101010001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0001000101110101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111000001001101001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011101001000001001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100100100001001001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111101101100101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010100011010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011001010010100001000000;
expected_data = 28'b1101101001000000000000000000;
@(next_data);

send_data = 28'b0000011001110001000010000000;
expected_data = 28'b0101001100000000000000000000;
@(next_data);

send_data = 28'b1000001101111110100011000000;
expected_data = 28'b0001101100000000000000000000;
@(next_data);

send_data = 28'b0000101000111000000100000000;
expected_data = 28'b0100000100000000000000000000;
@(next_data);

send_data = 28'b1001111101011100000101000000;
expected_data = 28'b0001010000000000000000000000;
@(next_data);

send_data = 28'b1001001100001101000110000000;
expected_data = 28'b1101000001000000000000000000;
@(next_data);

send_data = 28'b0101000001111000100111000000;
expected_data = 28'b1110110101000000000000000000;
@(next_data);

send_data = 28'b0110011001000000001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110001001111001001001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0101000000111111101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1100100001110111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111110100000101001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111001111000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000000100100010001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100011101110110101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011110001001001100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111101000001000001000000;
expected_data = 28'b1100111101000000000000000000;
@(next_data);

send_data = 28'b0010101101110010000010000000;
expected_data = 28'b1001110101000000000000000000;
@(next_data);

send_data = 28'b1010111000100101000011000000;
expected_data = 28'b0011000000000000000000000000;
@(next_data);

send_data = 28'b0100000001100111100100000000;
expected_data = 28'b0101011100000000000000000000;
@(next_data);

send_data = 28'b1010100100100100000101000000;
expected_data = 28'b1000000001100000000000000000;
@(next_data);

send_data = 28'b1101001001110011000110000000;
expected_data = 28'b1111110101000000000000000000;
@(next_data);

send_data = 28'b0101101100101111000111000000;
expected_data = 28'b1010111001000000000000000000;
@(next_data);

send_data = 28'b1100100001101000001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1101011000100001101001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1000111100111110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0111011101111101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111011100001011001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011110000011011101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110101111111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010101101011011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100000111101000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010111001111000100001000000;
expected_data = 28'b0000001000110000000000000000;
@(next_data);

send_data = 28'b1110011100100111000010000000;
expected_data = 28'b0101111100000000000000000000;
@(next_data);

send_data = 28'b0011010000011000000011000000;
expected_data = 28'b0101011000000000000000000000;
@(next_data);

send_data = 28'b1101001100000010000100000000;
expected_data = 28'b0001101000000000000000000000;
@(next_data);

send_data = 28'b1111111000111000100101000000;
expected_data = 28'b1010011001000000000000000000;
@(next_data);

send_data = 28'b1101111000001001000110000000;
expected_data = 28'b1000000101000000000000000000;
@(next_data);

send_data = 28'b0101010100001110000111000000;
expected_data = 28'b1010001001000000000000000000;
@(next_data);

send_data = 28'b0011101001001001101000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0010010001111000101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0111100001101011001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010101000011111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111001100111000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011110101100011101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111011000000110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101101000100011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011010101011110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111000000011001100001000000;
expected_data = 28'b1111000101000000000000000000;
@(next_data);

send_data = 28'b1011011101110101000010000000;
expected_data = 28'b1100001101000000000000000000;
@(next_data);

send_data = 28'b0010110100111111000011000000;
expected_data = 28'b1010001001000000000000000000;
@(next_data);

send_data = 28'b1100001001011111100100000000;
expected_data = 28'b0001011000000000000000000000;
@(next_data);

send_data = 28'b1011000100000001000101000000;
expected_data = 28'b1000010001000000000000000000;
@(next_data);

send_data = 28'b1110101100010010000110000000;
expected_data = 28'b1110100101000000000000000000;
@(next_data);

send_data = 28'b0111110000110010100111000000;
expected_data = 28'b1001010101000000000000000000;
@(next_data);

send_data = 28'b1101001000001011001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0110010000001010101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1011001101001001101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0000010000010100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101110001100010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101111001100100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001100101011001001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111001111011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100010000010001000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100101100011111000001000000;
expected_data = 28'b1110011001000000000000000000;
@(next_data);

send_data = 28'b0110111101111011100010000000;
expected_data = 28'b1111010101000000000000000000;
@(next_data);

send_data = 28'b1100100100011101100011000000;
expected_data = 28'b0110011100000000000000000000;
@(next_data);

send_data = 28'b1110010101010011100100000000;
expected_data = 28'b0110010000000000000000000000;
@(next_data);

send_data = 28'b0110111100111111000101000000;
expected_data = 28'b1100101001000000000000000000;
@(next_data);

send_data = 28'b1000001100001101100110000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b0010010101011000000111000000;
expected_data = 28'b1111110101000000000000000000;
@(next_data);

send_data = 28'b0111110101010000001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100100101000001101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0100001000011000001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0100001100101100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111010101011100101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001100000001111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010111001010100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101100000101100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110100110111100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011110001100001100001000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b0011101100011000000010000000;
expected_data = 28'b0111111100000000000000000000;
@(next_data);

send_data = 28'b0101000001010010100011000000;
expected_data = 28'b1111010001000000000000000000;
@(next_data);

send_data = 28'b1110110000101110100100000000;
expected_data = 28'b0010100000000000000000000000;
@(next_data);

send_data = 28'b0111101000010010000101000000;
expected_data = 28'b1101100001000000000000000000;
@(next_data);

send_data = 28'b1000100000110111000110000000;
expected_data = 28'b0100011100000000000000000000;
@(next_data);

send_data = 28'b1100000001010100000111000000;
expected_data = 28'b1111100001000000000000000000;
@(next_data);

send_data = 28'b0000001000110111001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001110001100011101001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b0111110101010000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0011101101010101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101101001110011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111101000110001101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100001100010010001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000010000011000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100010000101110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100100010100000001000000;
expected_data = 28'b0010000000110000000000000000;
@(next_data);

send_data = 28'b1010000001100010100010000000;
expected_data = 28'b1111000101000000000000000000;
@(next_data);

send_data = 28'b0010001000011001100011000000;
expected_data = 28'b1001101001000000000000000000;
@(next_data);

send_data = 28'b0101110100111100100100000000;
expected_data = 28'b0001000100000000000000000000;
@(next_data);

send_data = 28'b1010110001110101000101000000;
expected_data = 28'b1011101001000000000000000000;
@(next_data);

send_data = 28'b0011011000000110000110000000;
expected_data = 28'b1111101001000000000000000000;
@(next_data);

send_data = 28'b1101000100011001000111000000;
expected_data = 28'b0011011000000000000000000000;
@(next_data);

send_data = 28'b1111110101011011101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1011110100010010101001000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b0001010000101010001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0101011100010111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1000000001110010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010101101110010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011111001100111101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011001101000001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111001001001101100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100110101000110100001000000;
expected_data = 28'b0000110100010000000000000000;
@(next_data);

send_data = 28'b0111110000101111100010000000;
expected_data = 28'b0100000000100000000000000000;
@(next_data);

send_data = 28'b1011100101001001000011000000;
expected_data = 28'b1101110001000000000000000000;
@(next_data);

send_data = 28'b1001101001000101100100000000;
expected_data = 28'b0101110000000000000000000000;
@(next_data);

send_data = 28'b0111101000111110000101000000;
expected_data = 28'b0011010000000000000000000000;
@(next_data);

send_data = 28'b0001111000101110000110000000;
expected_data = 28'b0100011100000000000000000000;
@(next_data);

send_data = 28'b1111100100110101100111000000;
expected_data = 28'b0001111000000000000000000000;
@(next_data);

send_data = 28'b1110010101010011101000000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b1010011101001100001001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0001000100010110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0001101100011001101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1011000100011110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110100101011000001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101111001100110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000001000011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111100001101011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110000001100101000001000000;
expected_data = 28'b0100111100010000000000000000;
@(next_data);

send_data = 28'b0000001100001111100010000000;
expected_data = 28'b0010101000000000000000000000;
@(next_data);

send_data = 28'b1010001101010101000011000000;
expected_data = 28'b1110001101000000000000000000;
@(next_data);

send_data = 28'b1101100100001100100100000000;
expected_data = 28'b0101000100000000000000000000;
@(next_data);

send_data = 28'b1110111100100000000101000000;
expected_data = 28'b1011001001000000000000000000;
@(next_data);

send_data = 28'b0010110000011110100110000000;
expected_data = 28'b1001100001000000000000000000;
@(next_data);

send_data = 28'b1110110001010011000111000000;
expected_data = 28'b0010110000000000000000000000;
@(next_data);

send_data = 28'b0000011100110011001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110100101101001001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1101010101000101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010010100011011101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1001001000111001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110101000010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011101101011011001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101110101010110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000111101011000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110110100110110100001000000;
expected_data = 28'b0100000000110000000000000000;
@(next_data);

send_data = 28'b1100000101001111000010000000;
expected_data = 28'b1000000001100000000000000000;
@(next_data);

send_data = 28'b1000100101001100100011000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b0010101001010011000100000000;
expected_data = 28'b0100010000000000000000000000;
@(next_data);

send_data = 28'b1010111000101010000101000000;
expected_data = 28'b0101010000000000000000000000;
@(next_data);

send_data = 28'b1010001100000011000110000000;
expected_data = 28'b1111100101000000000000000000;
@(next_data);

send_data = 28'b0111100000111000000111000000;
expected_data = 28'b1101110101000000000000000000;
@(next_data);

send_data = 28'b1000100100001000101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010111000100000101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0001011100011111101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010100001111011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0001110100000001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000010101101110101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100001001010000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111001101001110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100101101100001100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110100101011111100001000000;
expected_data = 28'b0000111000010000000000000000;
@(next_data);

send_data = 28'b1001101101110110000010000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b0010101101011010100011000000;
expected_data = 28'b1000100001000000000000000000;
@(next_data);

send_data = 28'b0111010101010011100100000000;
expected_data = 28'b0001010100000000000000000000;
@(next_data);

send_data = 28'b1111000101000110100101000000;
expected_data = 28'b1110101001000000000000000000;
@(next_data);

send_data = 28'b0001110101000011000110000000;
expected_data = 28'b1000100101000000000000000000;
@(next_data);

send_data = 28'b1000010101000110100111000000;
expected_data = 28'b0001110100000000000000000000;
@(next_data);

send_data = 28'b0110100101011111101000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b1011011000000011001001000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1110100001001100101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1111000000110001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010100000110000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100101110101001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101100001100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100011000011011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010001001111100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110001101011111100001000000;
expected_data = 28'b1011001101000000000000000000;
@(next_data);

send_data = 28'b1100111001001001100010000000;
expected_data = 28'b1101110001000000000000000000;
@(next_data);

send_data = 28'b0110001001000110000011000000;
expected_data = 28'b1010001001000000000000000000;
@(next_data);

send_data = 28'b0111101001000111000100000000;
expected_data = 28'b0011000100000000000000000000;
@(next_data);

send_data = 28'b1000110100111100000101000000;
expected_data = 28'b1111010001000000000000000000;
@(next_data);

send_data = 28'b1000110000000001100110000000;
expected_data = 28'b1100101101000000000000000000;
@(next_data);

send_data = 28'b0001000001111101100111000000;
expected_data = 28'b1111010001000000000000000000;
@(next_data);

send_data = 28'b0111110000111110001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101101101111111001001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1011001000101111001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0110000101010011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101110101111101001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010011101001010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100010000001110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101111101001010001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110001100111100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111111100010010000001000000;
expected_data = 28'b1111101101000000000000000000;
@(next_data);

send_data = 28'b1110111001001010000010000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b0001111001110011000011000000;
expected_data = 28'b1000010101000000000000000000;
@(next_data);

send_data = 28'b1101000001100001000100000000;
expected_data = 28'b0000111100000000000000000000;
@(next_data);

send_data = 28'b1110101100101101100101000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b0011110000011110100110000000;
expected_data = 28'b1001111001000000000000000000;
@(next_data);

send_data = 28'b0011000001110110100111000000;
expected_data = 28'b0011110000000000000000000000;
@(next_data);

send_data = 28'b0111000000100111101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000111001011110001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0011010001100101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0111100100010010101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0100000000011000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010011100111111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101010000010100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110000000000011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110101101010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111101100101110100001000000;
expected_data = 28'b1000001001010000000000000000;
@(next_data);

send_data = 28'b1110100100110100000010000000;
expected_data = 28'b1010011001000000000000000000;
@(next_data);

send_data = 28'b0110011001100000000011000000;
expected_data = 28'b0111111000000000000000000000;
@(next_data);

send_data = 28'b1110011101010001100100000000;
expected_data = 28'b0011001100000000000000000000;
@(next_data);

send_data = 28'b0001000100011001100101000000;
expected_data = 28'b1100111001000000000000000000;
@(next_data);

send_data = 28'b1100111100110101100110000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b0001001001101000000111000000;
expected_data = 28'b1011000101000000000000000000;
@(next_data);

send_data = 28'b1100101000011011001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101011101000101101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1000100001001000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0100101000111100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010110100110001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100000000001101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011100100011001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000010100001001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100100010101000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101101001001100001000000;
expected_data = 28'b1011001101000000000000000000;
@(next_data);

send_data = 28'b0000001101111111100010000000;
expected_data = 28'b0011100000000000000000000000;
@(next_data);

send_data = 28'b0101101100101000100011000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b0000011101000101000100000000;
expected_data = 28'b0010110100000000000000000000;
@(next_data);

send_data = 28'b1001100001011011000101000000;
expected_data = 28'b0000111000000000000000000000;
@(next_data);

send_data = 28'b0100000000011101100110000000;
expected_data = 28'b1101010001000000000000000000;
@(next_data);

send_data = 28'b1111110000100100100111000000;
expected_data = 28'b0100000000100000000000000000;
@(next_data);

send_data = 28'b1110100100010011101000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0101100100110111101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0001111001110001001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0000000100111001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101011101110001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001001000011000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001101001010010001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001111000111110101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100000100001000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111110101010010000001000000;
expected_data = 28'b1100101001000000000000000000;
@(next_data);

send_data = 28'b1101100001100001100010000000;
expected_data = 28'b0101100100000000000000000000;
@(next_data);

send_data = 28'b0011010100000011100011000000;
expected_data = 28'b1110010001000000000000000000;
@(next_data);

send_data = 28'b0100111101100010100100000000;
expected_data = 28'b0001101000000000000000000000;
@(next_data);

send_data = 28'b1011010000101000100101000000;
expected_data = 28'b1001111001000000000000000000;
@(next_data);

send_data = 28'b1110000101101010100110000000;
expected_data = 28'b1110111001000000000000000000;
@(next_data);

send_data = 28'b0100111000011001100111000000;
expected_data = 28'b1001111101000000000000000000;
@(next_data);

send_data = 28'b0000001000001000001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1100110100010001101001000000;
expected_data = 28'b0000111000000000000000000000;
@(next_data);

send_data = 28'b1100000000110000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110001100001111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1100101101111110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110001101101001001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111011000101111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011000011110101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111001000010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011100010100100001000000;
expected_data = 28'b1101001101000000000000000000;
@(next_data);

send_data = 28'b0101110101001010000010000000;
expected_data = 28'b1101111001000000000000000000;
@(next_data);

send_data = 28'b0100010101000101000011000000;
expected_data = 28'b0011011000000000000000000000;
@(next_data);

send_data = 28'b1011011101001111000100000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b0011000000010101000101000000;
expected_data = 28'b0110111000000000000000000000;
@(next_data);

send_data = 28'b0101111001101011100110000000;
expected_data = 28'b0010100000000000000000000000;
@(next_data);

send_data = 28'b0111110101010001100111000000;
expected_data = 28'b0101111000000000000000000000;
@(next_data);

send_data = 28'b0010001101101011001000000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0000001100001101101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1000110100010101001010000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0100101101011111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0110101101111001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011001100110100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010010001011111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110111101000000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101001100101011000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011010000110111100001000000;
expected_data = 28'b1010100101000000000000000000;
@(next_data);

send_data = 28'b1110000001100101100010000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b1111001001011011000011000000;
expected_data = 28'b1101010001000000000000000000;
@(next_data);

send_data = 28'b0000111100101001100100000000;
expected_data = 28'b0111100100000000000000000000;
@(next_data);

send_data = 28'b0110111100001111000101000000;
expected_data = 28'b0001111000000000000000000000;
@(next_data);

send_data = 28'b1011100000101100000110000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b0001011101110011000111000000;
expected_data = 28'b1100100001000000000000000000;
@(next_data);

send_data = 28'b0011000100101100101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1110010101000001101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1111111001101010001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010110101100110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111010000000010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011000100010111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101001001001010101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100010001011010001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110100100000111100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110101101000000000001000000;
expected_data = 28'b1111100001000000000000000000;
@(next_data);

send_data = 28'b0000010000011101000010000000;
expected_data = 28'b0110101100000000000000000000;
@(next_data);

send_data = 28'b1011110101010010000011000000;
expected_data = 28'b1100000101000000000000000000;
@(next_data);

send_data = 28'b1111111000001110100100000000;
expected_data = 28'b0101111000000000000000000000;
@(next_data);

send_data = 28'b0110110101100001000101000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b0100101101110100000110000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b1100001101000000000111000000;
expected_data = 28'b0100101100000000000000000000;
@(next_data);

send_data = 28'b1110101000110110001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111010000011110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110010000110101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1001011101111110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111101000110001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010001100001010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011000010111101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100011000111010101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101100000000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110100000001101000001000000;
expected_data = 28'b0011110000000000000000000000;
@(next_data);

send_data = 28'b1100011000010100100010000000;
expected_data = 28'b1111001001000000000000000000;
@(next_data);

send_data = 28'b0011111001010000000011000000;
expected_data = 28'b0001000000100000000000000000;
@(next_data);

send_data = 28'b0000010000010110000100000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b1011110000110010000101000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1100101001000110100110000000;
expected_data = 28'b1110001001000000000000000000;
@(next_data);

send_data = 28'b0011111100010111000111000000;
expected_data = 28'b1011011001000000000000000000;
@(next_data);

send_data = 28'b1110010001101111101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0100100101110010001001000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0110100000111001001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010101100011100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110011100011110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110101001100010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010000100100111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100000001001110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100100100111011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001000101011010000001000000;
expected_data = 28'b1100000001000000000000000000;
@(next_data);

send_data = 28'b0111101100101100100010000000;
expected_data = 28'b0010010100000000000000000000;
@(next_data);

send_data = 28'b0010010100011001000011000000;
expected_data = 28'b1101110101000000000000000000;
@(next_data);

send_data = 28'b0111100101010100000100000000;
expected_data = 28'b0001001000000000000000000000;
@(next_data);

send_data = 28'b1000100000000100100101000000;
expected_data = 28'b1111001001000000000000000000;
@(next_data);

send_data = 28'b0011111001100011000110000000;
expected_data = 28'b1100110001000000000000000000;
@(next_data);

send_data = 28'b0110000001110001100111000000;
expected_data = 28'b0011111000000000000000000000;
@(next_data);

send_data = 28'b1000110000111100001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001010101100110101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0000101001110100001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010011101010000101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000000001011001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111110001001111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101011100010111101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001010100011101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110110101011001000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110001100111111100001000000;
expected_data = 28'b1001111101010000000000000000;
@(next_data);

send_data = 28'b1101000000000001100010000000;
expected_data = 28'b1001110001000000000000000000;
@(next_data);

send_data = 28'b0011101100001100000011000000;
expected_data = 28'b0010110000000000000000000000;
@(next_data);

send_data = 28'b1000110101011000000100000000;
expected_data = 28'b0001110100000000000000000000;
@(next_data);

send_data = 28'b1001010100111000000101000000;
expected_data = 28'b0001101000000000000000000000;
@(next_data);

send_data = 28'b0000101101000101000110000000;
expected_data = 28'b1101111101000000000000000000;
@(next_data);

send_data = 28'b0001011001100110100111000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0010100001111010001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0010001000000001101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1010001100100001101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0101111001001001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0110000001110001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110100101011111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011100101000001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011110101001100101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100101110110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111010000110000100001000000;
expected_data = 28'b1100011001010000000000000000;
@(next_data);

send_data = 28'b1100101001101100000010000000;
expected_data = 28'b0001010100000000000000000000;
@(next_data);

send_data = 28'b0101111100100100100011000000;
expected_data = 28'b1110110101000000000000000000;
@(next_data);

send_data = 28'b0100011100101110100100000000;
expected_data = 28'b0010111100000000000000000000;
@(next_data);

send_data = 28'b0011110000000110000101000000;
expected_data = 28'b1000111001000000000000000000;
@(next_data);

send_data = 28'b1110101100100100100110000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b0110010100101000000111000000;
expected_data = 28'b1001010101000000000000000000;
@(next_data);

send_data = 28'b1101011100000101001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101000100100101001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0110010000110110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011110101001110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111101101110000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101100001111010001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110000111010101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100110000011011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001011100101100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110111101111101000001000000;
expected_data = 28'b1111000001000000000000000000;
@(next_data);

send_data = 28'b1100010100000001000010000000;
expected_data = 28'b1001010101000000000000000000;
@(next_data);

send_data = 28'b1000100101111001000011000000;
expected_data = 28'b0011100000000000000000000000;
@(next_data);

send_data = 28'b1000011001011111100100000000;
expected_data = 28'b0100010000000000000000000000;
@(next_data);

send_data = 28'b0111001000000110000101000000;
expected_data = 28'b0000110000000000000000000000;
@(next_data);

send_data = 28'b1111000101110100000110000000;
expected_data = 28'b0100101100000000000000000000;
@(next_data);

send_data = 28'b0110111000000100000111000000;
expected_data = 28'b1000111101000000000000000000;
@(next_data);

send_data = 28'b1000110100110011001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001101100001110001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1101010101100110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1100011101000111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1001110101011100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100001100100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111000001010100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110101101100111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100000010000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001101101010001000001000000;
expected_data = 28'b1010100001000000000000000000;
@(next_data);

send_data = 28'b0111010100010000000010000000;
expected_data = 28'b0011100100000000000000000000;
@(next_data);

send_data = 28'b1100101100111101100011000000;
expected_data = 28'b1010101001000000000000000000;
@(next_data);

send_data = 28'b0000010001101110100100000000;
expected_data = 28'b0110010100000000000000000000;
@(next_data);

send_data = 28'b1100000100101010100101000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1000100001100011100110000000;
expected_data = 28'b1010000101000000000000000000;
@(next_data);

send_data = 28'b0110010101100101000111000000;
expected_data = 28'b1111100001000000000000000000;
@(next_data);

send_data = 28'b0001100001011000001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0001000101010110101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1101100000100000001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1001100100110011101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110101000110110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101000000111110101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001101100011100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101110100100111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110011100110010000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101010100110100000001000000;
expected_data = 28'b0100101100010000000000000000;
@(next_data);

send_data = 28'b1110100000100110000010000000;
expected_data = 28'b0011110100000000000000000000;
@(next_data);

send_data = 28'b0100101101000001000011000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b0100111001011011100100000000;
expected_data = 28'b0010010100000000000000000000;
@(next_data);

send_data = 28'b0100110101000010100101000000;
expected_data = 28'b1001110001000000000000000000;
@(next_data);

send_data = 28'b0111001001011110100110000000;
expected_data = 28'b0110101100000000000000000000;
@(next_data);

send_data = 28'b1001100001010001000111000000;
expected_data = 28'b0111001000000000000000000000;
@(next_data);

send_data = 28'b0001111001000011001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101110001110100101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1010010000001101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0110100000110000101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101110001111101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111100000110101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001101101011100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111110001101111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100010000011111100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001001000001001100001000000;
expected_data = 28'b0000001100010000000000000000;
@(next_data);

send_data = 28'b1000001000001011100010000000;
expected_data = 28'b1000000101000000000000000000;
@(next_data);

send_data = 28'b0100101101101110100011000000;
expected_data = 28'b0110101000000000000000000000;
@(next_data);

send_data = 28'b1100110100100011000100000000;
expected_data = 28'b0010010100000000000000000000;
@(next_data);

send_data = 28'b1101000101111000100101000000;
expected_data = 28'b1001101001000000000000000000;
@(next_data);

send_data = 28'b1100101000001100100110000000;
expected_data = 28'b1011100101000000000000000000;
@(next_data);

send_data = 28'b0110111101101010000111000000;
expected_data = 28'b1011011001000000000000000000;
@(next_data);

send_data = 28'b0001110000111110001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0011110100111001101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1100101100010100001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0111111101111000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0100100000101011001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111110000010100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011100000011001001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101001110001001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000100101100010000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101111100010001100001000000;
expected_data = 28'b1100110101000000000000000000;
@(next_data);

send_data = 28'b1111111101000101000010000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b0010001001001101000011000000;
expected_data = 28'b1000101001000000000000000000;
@(next_data);

send_data = 28'b1100000100111100100100000000;
expected_data = 28'b0001000100000000000000000000;
@(next_data);

send_data = 28'b1010000101010011000101000000;
expected_data = 28'b1000001001000000000000000000;
@(next_data);

send_data = 28'b0000001101010000100110000000;
expected_data = 28'b1111000101000000000000000000;
@(next_data);

send_data = 28'b0110011101101111000111000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b0110100100010000101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1000111101010011101001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b0011010101010111101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0100001001011111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101101000110101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100000011100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001000000010100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010001001110111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111100101111101100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110000101100111100001000000;
expected_data = 28'b0111010000010000000000000000;
@(next_data);

send_data = 28'b0111011000010010100010000000;
expected_data = 28'b1010111001000000000000000000;
@(next_data);

send_data = 28'b0100000000000000100011000000;
expected_data = 28'b1010110001000000000000000000;
@(next_data);

send_data = 28'b0100001000011100100100000000;
expected_data = 28'b0010000000100000000000000000;
@(next_data);

send_data = 28'b1010011000110101000101000000;
expected_data = 28'b1000010001000000000000000000;
@(next_data);

send_data = 28'b1110100001001011000110000000;
expected_data = 28'b1111010101000000000000000000;
@(next_data);

send_data = 28'b0001011100111001100111000000;
expected_data = 28'b1001100001000000000000000000;
@(next_data);

send_data = 28'b0011001001111101101000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b1100000101001011101001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0010001100110110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010111001010110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0001010100001110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111100000101111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001101001001100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101010101101011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110001110100000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101010100000011100001000000;
expected_data = 28'b1001010001010000000000000000;
@(next_data);

send_data = 28'b0101000101110001000010000000;
expected_data = 28'b1101001001000000000000000000;
@(next_data);

send_data = 28'b0010111101000111100011000000;
expected_data = 28'b0100110000000000000000000000;
@(next_data);

send_data = 28'b0011111000110010000100000000;
expected_data = 28'b0001011100000000000000000000;
@(next_data);

send_data = 28'b0110010101011101000101000000;
expected_data = 28'b0111110000000000000000000000;
@(next_data);

send_data = 28'b1001101001010110000110000000;
expected_data = 28'b0101011100000000000000000000;
@(next_data);

send_data = 28'b0010110001000000000111000000;
expected_data = 28'b1110011001000000000000000000;
@(next_data);

send_data = 28'b0111110101000100001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101110100001000001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0010110101001010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101011101101100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101010000100100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001110100111011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010001111001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000110101010001001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010101000001100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001000100111001000001000000;
expected_data = 28'b1001100001000000000000000000;
@(next_data);

send_data = 28'b0101011100011000100010000000;
expected_data = 28'b1110001101000000000000000000;
@(next_data);

send_data = 28'b1000110101111101100011000000;
expected_data = 28'b1001100101000000000000000000;
@(next_data);

send_data = 28'b0111111001101010000100000000;
expected_data = 28'b0100011000000000000000000000;
@(next_data);

send_data = 28'b1111100101100110000101000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b1001011000001010100110000000;
expected_data = 28'b1000010101000000000000000000;
@(next_data);

send_data = 28'b0110110100010100100111000000;
expected_data = 28'b1110101001000000000000000000;
@(next_data);

send_data = 28'b0010011000011111001000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1000010101001010101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0100010101101011001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110100101001000101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1100110101100000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101110100000111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101010100010001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001111001001000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111110101011111100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000001000110111100001000000;
expected_data = 28'b1011110001010000000000000000;
@(next_data);

send_data = 28'b1010001101111110000010000000;
expected_data = 28'b1110110101000000000000000000;
@(next_data);

send_data = 28'b0001010000011010000011000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b1010000100101011100100000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b0001010001000110100101000000;
expected_data = 28'b0100001000000000000000000000;
@(next_data);

send_data = 28'b1010110100111010100110000000;
expected_data = 28'b0001111000000000000000000000;
@(next_data);

send_data = 28'b1011011101100101100111000000;
expected_data = 28'b1101001101000000000000000000;
@(next_data);

send_data = 28'b1110010101000101101000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b1111000000110000101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1011001000101010001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010100100110001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1000100100101001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011011100111000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110001000110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111000100001101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011001000011000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110100001011100001000000;
expected_data = 28'b0000110000010000000000000000;
@(next_data);

send_data = 28'b1010101001010010000010000000;
expected_data = 28'b0011101000000000000000000000;
@(next_data);

send_data = 28'b1001001100101111100011000000;
expected_data = 28'b1111000101000000000000000000;
@(next_data);

send_data = 28'b0001111101011011100100000000;
expected_data = 28'b0100100100000000000000000000;
@(next_data);

send_data = 28'b0000001101010001000101000000;
expected_data = 28'b0011111000000000000000000000;
@(next_data);

send_data = 28'b0000101001110111000110000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0000001001111101000111000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b0100011101101010001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1111001000110100001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0001011001010101101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0111000100000111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0110110101100000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100001101010000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000000000100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011101111001001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101001011101000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011000000011011100001000000;
expected_data = 28'b0110010000010000000000000000;
@(next_data);

send_data = 28'b0011100100000000000010000000;
expected_data = 28'b1000011101000000000000000000;
@(next_data);

send_data = 28'b1111001101101110000011000000;
expected_data = 28'b1100011001000000000000000000;
@(next_data);

send_data = 28'b0100100001011001100100000000;
expected_data = 28'b0111100100000000000000000000;
@(next_data);

send_data = 28'b1010100000110101000101000000;
expected_data = 28'b1001000001000000000000000000;
@(next_data);

send_data = 28'b0011000000001010000110000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b0101110001000001100111000000;
expected_data = 28'b0011000000000000000000000000;
@(next_data);

send_data = 28'b1011000100111100101000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1111001000101010101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0110101001111000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011100001001000101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1011010101100011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010111100101011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111101110110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111110101111111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101000011010000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011111000101100100001000000;
expected_data = 28'b0110111000000000000000000000;
@(next_data);

send_data = 28'b0111010100110001100010000000;
expected_data = 28'b1110011101000000000000000000;
@(next_data);

send_data = 28'b0011001100100000000011000000;
expected_data = 28'b1110100101000000000000000000;
@(next_data);

send_data = 28'b0100010000000001000100000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b0111111001111100100101000000;
expected_data = 28'b1000100001000000000000000000;
@(next_data);

send_data = 28'b1111101001111100000110000000;
expected_data = 28'b0100000100000000000000000000;
@(next_data);

send_data = 28'b1110100100110101000111000000;
expected_data = 28'b1000011001000000000000000000;
@(next_data);

send_data = 28'b0110000101100110101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1111001101000101101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1111110101011001101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0000100000001110001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111010000001101001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100010000000001101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011000000000001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000001100101111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110000001100011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010011101011101100001000000;
expected_data = 28'b1010011101010000000000000000;
@(next_data);

send_data = 28'b1101101001001011000010000000;
expected_data = 28'b0001110000000000000000000000;
@(next_data);

send_data = 28'b0110110000101101100011000000;
expected_data = 28'b1011001101000000000000000000;
@(next_data);

send_data = 28'b0001000100101010100100000000;
expected_data = 28'b0011011000000000000000000000;
@(next_data);

send_data = 28'b1001100100001110100101000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b1001100100010000000110000000;
expected_data = 28'b1101010101000000000000000000;
@(next_data);

send_data = 28'b1110101001110101100111000000;
expected_data = 28'b1110011101000000000000000000;
@(next_data);

send_data = 28'b0110110100010000101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1000110000010011001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0111100101111011001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1000011000001100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1001011000110011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110000001101000001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111001001000110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110001100110111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001110100011110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111000101010100001000000;
expected_data = 28'b0101100100000000000000000000;
@(next_data);

send_data = 28'b0011111001101100000010000000;
expected_data = 28'b0001101100000000000000000000;
@(next_data);

send_data = 28'b1100111100011001000011000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b1000100100101010000100000000;
expected_data = 28'b0110011100000000000000000000;
@(next_data);

send_data = 28'b1010010000101110000101000000;
expected_data = 28'b0001001000000000000000000000;
@(next_data);

send_data = 28'b1001101001000101100110000000;
expected_data = 28'b1111011001000000000000000000;
@(next_data);

send_data = 28'b1011001100111101100111000000;
expected_data = 28'b1110011001000000000000000000;
@(next_data);

send_data = 28'b1100001001011100001000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1111000001111101001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1101111100011011101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0110111100010101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101111000101000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111101101001111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111101000100011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000101011101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100110000101010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011000101101011000001000000;
expected_data = 28'b1010000101000000000000000000;
@(next_data);

send_data = 28'b1100110001110010000010000000;
expected_data = 28'b1110011101000000000000000000;
@(next_data);

send_data = 28'b1010001000000010000011000000;
expected_data = 28'b1101011101000000000000000000;
@(next_data);

send_data = 28'b0101101001001111100100000000;
expected_data = 28'b0101000100000000000000000000;
@(next_data);

send_data = 28'b1110001001111001000101000000;
expected_data = 28'b1011010001000000000000000000;
@(next_data);

send_data = 28'b1101111101011000100110000000;
expected_data = 28'b1001001101000000000000000000;
@(next_data);

send_data = 28'b1011010001100011100111000000;
expected_data = 28'b1010000101000000000000000000;
@(next_data);

send_data = 28'b0010011001101001001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1110011101001001001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1000011100110101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0001011000010101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110100100111001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010001100000100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101100100110001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101011000000111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001110101100110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110010101010010100001000000;
expected_data = 28'b0110101000010000000000000000;
@(next_data);

send_data = 28'b0000100101110101000010000000;
expected_data = 28'b1100000001000000000000000000;
@(next_data);

send_data = 28'b0100011100100100000011000000;
expected_data = 28'b0001110000000000000000000000;
@(next_data);

send_data = 28'b0000110001100110100100000000;
expected_data = 28'b0010001100000000000000000000;
@(next_data);

send_data = 28'b0010111001101010100101000000;
expected_data = 28'b0001100000000000000000000000;
@(next_data);

send_data = 28'b1010000100111111100110000000;
expected_data = 28'b0011100100000000000000000000;
@(next_data);

send_data = 28'b0111001001011001100111000000;
expected_data = 28'b1101111101000000000000000000;
@(next_data);

send_data = 28'b0011100001010010101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1101001100011000101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0010000101111110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110011100010110001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010101000110000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000000000110000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111010001000110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111010000110100101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001110000101011000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001011101110001100001000000;
expected_data = 28'b0111001000000000000000000000;
@(next_data);

send_data = 28'b1101001001001001000010000000;
expected_data = 28'b0111010000000000000000000000;
@(next_data);

send_data = 28'b0011011001010101100011000000;
expected_data = 28'b1011111101000000000000000000;
@(next_data);

send_data = 28'b1111111000110111100100000000;
expected_data = 28'b0001101100000000000000000000;
@(next_data);

send_data = 28'b1111110001011001100101000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b0111010100101111000110000000;
expected_data = 28'b1000001001000000000000000000;
@(next_data);

send_data = 28'b1000101100101101100111000000;
expected_data = 28'b0111010100000000000000000000;
@(next_data);

send_data = 28'b0110110000101111001000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1010111001101001101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1011011101101001101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0110011100111101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110110101010100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101000001010111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000101101110100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011000000001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100001001100000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000110100110011000001000000;
expected_data = 28'b0100000000110000000000000000;
@(next_data);

send_data = 28'b0101110001111111100010000000;
expected_data = 28'b0110101100000000000000000000;
@(next_data);

send_data = 28'b1111111100001010100011000000;
expected_data = 28'b0101110000000000000000000000;
@(next_data);

send_data = 28'b0110101000000110000100000000;
expected_data = 28'b0111111100000000000000000000;
@(next_data);

send_data = 28'b0101011001111000100101000000;
expected_data = 28'b1101010001000000000000000000;
@(next_data);

send_data = 28'b0100010000010101100110000000;
expected_data = 28'b0111110100000000000000000000;
@(next_data);

send_data = 28'b1011011000001001100111000000;
expected_data = 28'b0100010000000000000000000000;
@(next_data);

send_data = 28'b0001000000010001001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0000011100010101101001000000;
expected_data = 28'b0000110100000000000000000000;
@(next_data);

send_data = 28'b1010100000100110001010000000;
expected_data = 28'b0111111100000000000000000000;
@(next_data);

send_data = 28'b0011001001001100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101010101100101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110110001011010001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011010000000111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100111000100110101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111110100011011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010001011111000001000000;
expected_data = 28'b0011010000010000000000000000;
@(next_data);

send_data = 28'b0011010001100100000010000000;
expected_data = 28'b0001101000000000000000000000;
@(next_data);

send_data = 28'b0100100101010010000011000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b0101110100010010100100000000;
expected_data = 28'b0010010000000000000000000000;
@(next_data);

send_data = 28'b1101111101010110100101000000;
expected_data = 28'b1011101001000000000000000000;
@(next_data);

send_data = 28'b0101001000011111000110000000;
expected_data = 28'b1011000001000000000000000000;
@(next_data);

send_data = 28'b1100000100110100100111000000;
expected_data = 28'b0101001000000000000000000000;
@(next_data);

send_data = 28'b0100101000001001001000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b0000100001010010101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1010111100011101001010000000;
expected_data = 28'b1111111111000000000000000000;
@(next_data);

send_data = 28'b1111110100011111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101111000100011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100001101110101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101110100001001001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010010101111000001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110001100110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101000100011001000001000000;
expected_data = 28'b0111100000010000000000000000;
@(next_data);

send_data = 28'b0011111000000000000010000000;
expected_data = 28'b1110001101000000000000000000;
@(next_data);

send_data = 28'b1101011001010111000011000000;
expected_data = 28'b1100000101000000000000000000;
@(next_data);

send_data = 28'b1100000100011000100100000000;
expected_data = 28'b0110101100000000000000000000;
@(next_data);

send_data = 28'b1101010001011101100101000000;
expected_data = 28'b1000001001000000000000000000;
@(next_data);

send_data = 28'b0011100100110011000110000000;
expected_data = 28'b1011111001000000000000000000;
@(next_data);

send_data = 28'b1001001000010000000111000000;
expected_data = 28'b0011100100000000000000000000;
@(next_data);

send_data = 28'b0001011100100000101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111001100110001101001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1101101101110110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1001001000101111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101110001001000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101101000010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111000111111101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111101100101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111001110100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010000001100001000001000000;
expected_data = 28'b0000011100010000000000000000;
@(next_data);

send_data = 28'b1011011100010111000010000000;
expected_data = 28'b0110001000000000000000000000;
@(next_data);

send_data = 28'b0111111001100000100011000000;
expected_data = 28'b0110011000000000000000000000;
@(next_data);

send_data = 28'b0101010001010000000100000000;
expected_data = 28'b0011111100000000000000000000;
@(next_data);

send_data = 28'b0000011101010101000101000000;
expected_data = 28'b1010100001000000000000000000;
@(next_data);

send_data = 28'b1110110001110101000110000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0010011100011010100111000000;
expected_data = 28'b1001010001000000000000000000;
@(next_data);

send_data = 28'b0100111001011111001000000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b1010000100100001101001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1001010100010011101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101011100010011101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111101100001000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101001100110101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010100101100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110010101111100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001010100001100000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011100000010010100001000000;
expected_data = 28'b1010110101000000000000000000;
@(next_data);

send_data = 28'b0011001100101001100010000000;
expected_data = 28'b1001110101000000000000000000;
@(next_data);

send_data = 28'b0011000001010010100011000000;
expected_data = 28'b1001111101000000000000000000;
@(next_data);

send_data = 28'b1010111101101101100100000000;
expected_data = 28'b0001100000000000000000000000;
@(next_data);

send_data = 28'b1110001101011111100101000000;
expected_data = 28'b0101111000000000000000000000;
@(next_data);

send_data = 28'b1011010101000100000110000000;
expected_data = 28'b1001001001000000000000000000;
@(next_data);

send_data = 28'b1001011001101110100111000000;
expected_data = 28'b1100101101000000000000000000;
@(next_data);

send_data = 28'b1001110001000111101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1000001101101011001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1001111100010011001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1100100001111011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1011110100010110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110010000011111001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101100100001100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111100101100011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010101101101101100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101011001100101100001000000;
expected_data = 28'b0000011000010000000000000000;
@(next_data);

send_data = 28'b1001111101110100100010000000;
expected_data = 28'b1001110101000000000000000000;
@(next_data);

send_data = 28'b1111010100101011100011000000;
expected_data = 28'b1000100101000000000000000000;
@(next_data);

send_data = 28'b0100000000100000100100000000;
expected_data = 28'b0111101000000000000000000000;
@(next_data);

send_data = 28'b0110110001111011100101000000;
expected_data = 28'b1000000001100000000000000000;
@(next_data);

send_data = 28'b0011011100111100000110000000;
expected_data = 28'b0101101000000000000000000000;
@(next_data);

send_data = 28'b0000111001000010000111000000;
expected_data = 28'b0011011100000000000000000000;
@(next_data);

send_data = 28'b1000011001011001001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010000100110100001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0000111101001111101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0111100100110100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111111100100000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101100101100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011100001011010001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111011101011111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101000101010110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111001101101100001000000;
expected_data = 28'b0111110100010000000000000000;
@(next_data);

send_data = 28'b0100000001110000100010000000;
expected_data = 28'b1001010101000000000000000000;
@(next_data);

send_data = 28'b1110110000000111000011000000;
expected_data = 28'b0101111000000000000000000000;
@(next_data);

send_data = 28'b0101000000010100100100000000;
expected_data = 28'b0111011000000000000000000000;
@(next_data);

send_data = 28'b0011110000000100000101000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b0110110100110100000110000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b1101010101100111000111000000;
expected_data = 28'b0110110100000000000000000000;
@(next_data);

send_data = 28'b0110101100001110101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0001111001111111001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0101100001100000001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0001011000101000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111010101010001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010000101100101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110101001001010001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010111101010000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101001001111110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000111000011010100001000000;
expected_data = 28'b0100111000010000000000000000;
@(next_data);

send_data = 28'b1011001101010010000010000000;
expected_data = 28'b0011101100000000000000000000;
@(next_data);

send_data = 28'b0100111100011100100011000000;
expected_data = 28'b1110100001000000000000000000;
@(next_data);

send_data = 28'b1111111101110010100100000000;
expected_data = 28'b0010011100000000000000000000;
@(next_data);

send_data = 28'b1000011100101111100101000000;
expected_data = 28'b1111111001000000000000000000;
@(next_data);

send_data = 28'b1010101001000000000110000000;
expected_data = 28'b1100010001000000000000000000;
@(next_data);

send_data = 28'b0100100101001100000111000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b1000000001011111001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011001000101000101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0100001000010110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110001101011011101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010101001001101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011010100101111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110110001001110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000110000110011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111000011011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001101100111000000001000000;
expected_data = 28'b1000010101000000000000000000;
@(next_data);

send_data = 28'b1110110000001000100010000000;
expected_data = 28'b1110101101000000000000000000;
@(next_data);

send_data = 28'b0110111000111110100011000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0100001101011110000100000000;
expected_data = 28'b0011011100000000000000000000;
@(next_data);

send_data = 28'b0001100100010001000101000000;
expected_data = 28'b1000011001000000000000000000;
@(next_data);

send_data = 28'b1001011100101111000110000000;
expected_data = 28'b0001010100000000000000000000;
@(next_data);

send_data = 28'b1110000001111011000111000000;
expected_data = 28'b1110100101000000000000000000;
@(next_data);

send_data = 28'b1101001000111101001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010111101101011101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110111000000001001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0011110101110000101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000001000111000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110101001011101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011000010011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001000000100000001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100000001011110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001001001101101100001000000;
expected_data = 28'b1111110101000000000000000000;
@(next_data);

send_data = 28'b0011100001000010000010000000;
expected_data = 28'b0100100100000000000000000000;
@(next_data);

send_data = 28'b1010111101011101000011000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b1110110101110111000100000000;
expected_data = 28'b0101011100000000000000000000;
@(next_data);

send_data = 28'b0101001100010110100101000000;
expected_data = 28'b1101101001000000000000000000;
@(next_data);

send_data = 28'b0011100100001101000110000000;
expected_data = 28'b0111101000000000000000000000;
@(next_data);

send_data = 28'b0010100000011010000111000000;
expected_data = 28'b0011100100000000000000000000;
@(next_data);

send_data = 28'b0100100000011000101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111001011100101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1101010001101010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1001011100100011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1011100100101110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011100101010110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011000000011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101011001001010101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111100101110100000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010100000111110100001000000;
expected_data = 28'b0110000100010000000000000000;
@(next_data);

send_data = 28'b0011110001100101100010000000;
expected_data = 28'b0101010100000000000000000000;
@(next_data);

send_data = 28'b1001010100000011000011000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1010010101011001100100000000;
expected_data = 28'b0100101000000000000000000000;
@(next_data);

send_data = 28'b0011001000001011100101000000;
expected_data = 28'b0100101000000000000000000000;
@(next_data);

send_data = 28'b1110100100100001000110000000;
expected_data = 28'b0010101100000000000000000000;
@(next_data);

send_data = 28'b1100100001101100000111000000;
expected_data = 28'b1001011101000000000000000000;
@(next_data);

send_data = 28'b1001111101011011001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010000001101110001001000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1100010001011001101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0111111001001101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110000101001011001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010000001000111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111001101000100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000111100000011001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010010000000110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110000001100000001000000;
expected_data = 28'b0011000000000000000000000000;
@(next_data);

send_data = 28'b1111010000011000100010000000;
expected_data = 28'b0011010000000000000000000000;
@(next_data);

send_data = 28'b1011011001010111000011000000;
expected_data = 28'b0011101000000000000000000000;
@(next_data);

send_data = 28'b1110101000011101000100000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b0100100100010110100101000000;
expected_data = 28'b1101010001000000000000000000;
@(next_data);

send_data = 28'b0101101101101110100110000000;
expected_data = 28'b0110110100000000000000000000;
@(next_data);

send_data = 28'b0111111001001110100111000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b0110110101101100101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0010111001101110001001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1110100100010000001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1001011001100100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110100000100011001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100000101110100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110000110110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011100110110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100000100111000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000000010000000001000000;
expected_data = 28'b1011000101000000000000000000;
@(next_data);

send_data = 28'b1011010100111011000010000000;
expected_data = 28'b0010000000100000000000000000;
@(next_data);

send_data = 28'b1100010000011101000011000000;
expected_data = 28'b0011110000000000000000000000;
@(next_data);

send_data = 28'b0001001101010110000100000000;
expected_data = 28'b0110001000000000000000000000;
@(next_data);

send_data = 28'b1100001100111010100101000000;
expected_data = 28'b0010011000000000000000000000;
@(next_data);

send_data = 28'b1001100000110101100110000000;
expected_data = 28'b1010001001000000000000000000;
@(next_data);

send_data = 28'b0001111100111100000111000000;
expected_data = 28'b1110100001000000000000000000;
@(next_data);

send_data = 28'b0001111100110000001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100100000101001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1100001000001101101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1001101101111001101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0001000001001001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001001100001110101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011001111000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001111001101100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101000101100000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010001100100000001000000;
expected_data = 28'b0000001000110000000000000000;
@(next_data);

send_data = 28'b0010110001101001100010000000;
expected_data = 28'b0110110000000000000000000000;
@(next_data);

send_data = 28'b1000011000110100100011000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101000100010100100100000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b0110001001010101100101000000;
expected_data = 28'b1010001001000000000000000000;
@(next_data);

send_data = 28'b0000010001110000100110000000;
expected_data = 28'b0101001100000000000000000000;
@(next_data);

send_data = 28'b1001101101001011000111000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1111110000000100001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0110101100111010001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0010100000001011101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0110001000111001101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111011001001011001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010011100100001101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010001001100011001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111101001000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000101111111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110001111010000001000000;
expected_data = 28'b0000111100010000000000000000;
@(next_data);

send_data = 28'b0101110101111100100010000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b1101110000010111100011000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b1010110001100100100100000000;
expected_data = 28'b0110111000000000000000000000;
@(next_data);

send_data = 28'b1000001100100010100101000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b0101100101011000000110000000;
expected_data = 28'b1100001001000000000000000000;
@(next_data);

send_data = 28'b1111011100101101000111000000;
expected_data = 28'b0101100100000000000000000000;
@(next_data);

send_data = 28'b0010000001000100001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1100010001101101101001000000;
expected_data = 28'b0000110100000000000000000000;
@(next_data);

send_data = 28'b0100101100000000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101011001101110001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000110100110010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010001000010110101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011000001011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110100001100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000001001001100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100011000100011000001000000;
expected_data = 28'b1001001101000000000000000000;
@(next_data);

send_data = 28'b1010010100001000100010000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011111101011110100011000000;
expected_data = 28'b0100101100000000000000000000;
@(next_data);

send_data = 28'b0000001001001101100100000000;
expected_data = 28'b0101111100000000000000000000;
@(next_data);

send_data = 28'b0001100000111000100101000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1010101101011110100110000000;
expected_data = 28'b0001010000000000000000000000;
@(next_data);

send_data = 28'b0101000100110001000111000000;
expected_data = 28'b1101010101000000000000000000;
@(next_data);

send_data = 28'b1000001001000110001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0101111101011110101001000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b1011010100011111101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1111110001111100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1010000000000110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100010000110010001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011000001000100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110001000010010101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100000100000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011011000001010000001000000;
expected_data = 28'b0001100100010000000000000000;
@(next_data);

send_data = 28'b1011100101011110000010000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b0011111100111100000011000000;
expected_data = 28'b1111101001000000000000000000;
@(next_data);

send_data = 28'b0000101101010011100100000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b1010110000001010000101000000;
expected_data = 28'b0001011000000000000000000000;
@(next_data);

send_data = 28'b0110001100110100100110000000;
expected_data = 28'b1111101001000000000000000000;
@(next_data);

send_data = 28'b1110000001000000100111000000;
expected_data = 28'b0110001100000000000000000000;
@(next_data);

send_data = 28'b1110111101011110001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100101100100110001001000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0100011001010110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1111000001100101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101010001000111001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110010000010101001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011000011010001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010111101010101001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101001100010101000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100100110111000001000000;
expected_data = 28'b1111110101000000000000000000;
@(next_data);

send_data = 28'b1010011000001001000010000000;
expected_data = 28'b1011011101000000000000000000;
@(next_data);

send_data = 28'b1000010001111111100011000000;
expected_data = 28'b0100101100000000000000000000;
@(next_data);

send_data = 28'b0101100001110111000100000000;
expected_data = 28'b0100001000000000000000000000;
@(next_data);

send_data = 28'b0110010001100110000101000000;
expected_data = 28'b1011000001000000000000000000;
@(next_data);

send_data = 28'b0100010001000100100110000000;
expected_data = 28'b0101011000000000000000000000;
@(next_data);

send_data = 28'b1111001001100010100111000000;
expected_data = 28'b0100010000000000000000000000;
@(next_data);

send_data = 28'b0000110101011010101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0011001100111001101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0011011101010000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110011001000101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010010001110100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111000100111100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100101010110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110111101100110101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000001100110100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010011000001110000001000000;
expected_data = 28'b0110110000000000000000000000;
@(next_data);

send_data = 28'b1101000001010011000010000000;
expected_data = 28'b0011101000000000000000000000;
@(next_data);

send_data = 28'b1100111100010100000011000000;
expected_data = 28'b1000100101000000000000000000;
@(next_data);

send_data = 28'b0101000000110100000100000000;
expected_data = 28'b0110011100000000000000000000;
@(next_data);

send_data = 28'b1111100101110110100101000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b0110100100110110100110000000;
expected_data = 28'b1000010101000000000000000000;
@(next_data);

send_data = 28'b1110110100111000100111000000;
expected_data = 28'b0110100100000000000000000000;
@(next_data);

send_data = 28'b0101100100000111001000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0101100001101011001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0001100101110011101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010101001010111101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110001100000110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111001100000000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111001111111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010001111000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101001000000111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100001001110000001000000;
expected_data = 28'b0110000000000000000000000000;
@(next_data);

send_data = 28'b1111001100111111100010000000;
expected_data = 28'b0011010000000000000000000000;
@(next_data);

send_data = 28'b0111011000000000100011000000;
expected_data = 28'b0111001100000000000000000000;
@(next_data);

send_data = 28'b0011001000000001100100000000;
expected_data = 28'b0011101100000000000000000000;
@(next_data);

send_data = 28'b1100000001000011000101000000;
expected_data = 28'b0110010000000000000000000000;
@(next_data);

send_data = 28'b0100011001101110000110000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b0100111100000001000111000000;
expected_data = 28'b0100011000000000000000000000;
@(next_data);

send_data = 28'b0010101000101001101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1001001001101000101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1101001101100010001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010000101110000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0011111001110100101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000100100010110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000010001010101001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100101010110101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000000000010010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011000010011000001000000;
expected_data = 28'b1010010101000000000000000000;
@(next_data);

send_data = 28'b0010010100001111100010000000;
expected_data = 28'b1010000001000000000000000000;
@(next_data);

send_data = 28'b1110101101101001000011000000;
expected_data = 28'b1100010101000000000000000000;
@(next_data);

send_data = 28'b0001011101010100100100000000;
expected_data = 28'b0111010100000000000000000000;
@(next_data);

send_data = 28'b1010001100101110000101000000;
expected_data = 28'b0010111000000000000000000000;
@(next_data);

send_data = 28'b1010001100001010000110000000;
expected_data = 28'b1111001001000000000000000000;
@(next_data);

send_data = 28'b1010111000010110100111000000;
expected_data = 28'b1101110101000000000000000000;
@(next_data);

send_data = 28'b1010110100000101101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0101001100111011101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1010100001111010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0100011100000000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0011100100110000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110101000001101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001001001010110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100111101101000101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010100001010111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111110101010101100001000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b1101001000111111100010000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b1011011000001100000011000000;
expected_data = 28'b0101001000000000000000000000;
@(next_data);

send_data = 28'b1110111000011100100100000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b0010010101110110000101000000;
expected_data = 28'b1101110001000000000000000000;
@(next_data);

send_data = 28'b1010010101100110100110000000;
expected_data = 28'b0011011100000000000000000000;
@(next_data);

send_data = 28'b1011100101101110100111000000;
expected_data = 28'b1101101101000000000000000000;
@(next_data);

send_data = 28'b1110011101011010001000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1010010001001001101001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0010111101010111101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010111100010101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1010111000100111101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110010001010100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011000111100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100000000110011101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011110001010010000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110000101101000000001000000;
expected_data = 28'b0110000000010000000000000000;
@(next_data);

send_data = 28'b1011111100000111100010000000;
expected_data = 28'b0011000100000000000000000000;
@(next_data);

send_data = 28'b0111100001000101100011000000;
expected_data = 28'b0100111100000000000000000000;
@(next_data);

send_data = 28'b0111111001000101100100000000;
expected_data = 28'b0011110000000000000000000000;
@(next_data);

send_data = 28'b0110001000110110000101000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b1100011000011011000110000000;
expected_data = 28'b0101001100000000000000000000;
@(next_data);

send_data = 28'b0011011000011100000111000000;
expected_data = 28'b1011101001000000000000000000;
@(next_data);

send_data = 28'b1011011101100010001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010011001010100101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0101100101010000001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1000011101011000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101000101000100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110000000110011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100001111011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101000001010111001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000010101111100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001111101111011000001000000;
expected_data = 28'b0111111000010000000000000000;
@(next_data);

send_data = 28'b0000100101011100100010000000;
expected_data = 28'b0110100100000000000000000000;
@(next_data);

send_data = 28'b1110011100001011100011000000;
expected_data = 28'b0100111100000000000000000000;
@(next_data);

send_data = 28'b0110100000110111100100000000;
expected_data = 28'b0111001100000000000000000000;
@(next_data);

send_data = 28'b0000110101100100000101000000;
expected_data = 28'b1101000001000000000000000000;
@(next_data);

send_data = 28'b1101100001111010100110000000;
expected_data = 28'b0000101100000000000000000000;
@(next_data);

send_data = 28'b0000001101001100100111000000;
expected_data = 28'b1010100001000000000000000000;
@(next_data);

send_data = 28'b1101001001010100101000000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b0001001101111010101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0111000001110101101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0001001000001110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1010111101101100101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101110101001110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011010101000111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110100000001111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010101001011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011111000011001100001000000;
expected_data = 28'b0011110000010000000000000000;
@(next_data);

send_data = 28'b0010010001101110100010000000;
expected_data = 28'b0000110100000000000000000000;
@(next_data);

send_data = 28'b1101010001110010100011000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0010001001010110100100000000;
expected_data = 28'b0110101000000000000000000000;
@(next_data);

send_data = 28'b0111000101010100000101000000;
expected_data = 28'b0100010000000000000000000000;
@(next_data);

send_data = 28'b0000011000010100100110000000;
expected_data = 28'b0100100100000000000000000000;
@(next_data);

send_data = 28'b0001011001001011000111000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1100010101100100001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0011101100110100101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0001001000010111001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010110000011001101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010101100000010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111000100100110101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110010100001011001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000100100110101001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011000110000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101000101100100001000000;
expected_data = 28'b0111011000000000000000000000;
@(next_data);

send_data = 28'b1101110100101010100010000000;
expected_data = 28'b1000001101000000000000000000;
@(next_data);

send_data = 28'b0010100000101000100011000000;
expected_data = 28'b0111011100000000000000000000;
@(next_data);

send_data = 28'b1111111000000011000100000000;
expected_data = 28'b0001010000000000000000000000;
@(next_data);

send_data = 28'b0111000100110011100101000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b1101001100110101000110000000;
expected_data = 28'b0100100100000000000000000000;
@(next_data);

send_data = 28'b0111110101111101100111000000;
expected_data = 28'b1010110101000000000000000000;
@(next_data);

send_data = 28'b1111011101000000001000000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0000100001011000101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0011101100111111001010000000;
expected_data = 28'b1111111111000000000000000000;
@(next_data);

send_data = 28'b0100101001110110001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000000001100011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100110000011000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011001110001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101000000111100101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100100010110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010100101110110100001000000;
expected_data = 28'b1101011001000000000000000000;
@(next_data);

send_data = 28'b0101100000111000000010000000;
expected_data = 28'b1100010001000000000000000000;
@(next_data);

send_data = 28'b1110001101111010000011000000;
expected_data = 28'b1101011101000000000000000000;
@(next_data);

send_data = 28'b0010001000010111100100000000;
expected_data = 28'b0111000100000000000000000000;
@(next_data);

send_data = 28'b1000100100001110000101000000;
expected_data = 28'b0100010000000000000000000000;
@(next_data);

send_data = 28'b0001101001100011000110000000;
expected_data = 28'b1100110101000000000000000000;
@(next_data);

send_data = 28'b0101111101100101100111000000;
expected_data = 28'b0001101000000000000000000000;
@(next_data);

send_data = 28'b1010010100010011101000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b0111101100011000101001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b0011100100110100001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1111100000111110001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0100001001101010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011010101011101001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100111101100000001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110110100110101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011101101000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111011100010111100001000000;
expected_data = 28'b1101100001000000000000000000;
@(next_data);

send_data = 28'b0001001101111101000010000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b0001110101001101100011000000;
expected_data = 28'b0001011000000000000000000000;
@(next_data);

send_data = 28'b1000111001101101100100000000;
expected_data = 28'b0000111000000000000000000000;
@(next_data);

send_data = 28'b1100101101001010000101000000;
expected_data = 28'b0001110000000000000000000000;
@(next_data);

send_data = 28'b0000110101100010000110000000;
expected_data = 28'b1010111001000000000000000000;
@(next_data);

send_data = 28'b1111101000100010000111000000;
expected_data = 28'b0000110100000000000000000000;
@(next_data);

send_data = 28'b1110010100000101001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110100000010001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1011010101111000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101101000100101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101111001101100101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000110000001001001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110111101110111101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101001001100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011010000001010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101000001011100001000000;
expected_data = 28'b1100100101000000000000000000;
@(next_data);

send_data = 28'b1110001000011000100010000000;
expected_data = 28'b1011110101000000000000000000;
@(next_data);

send_data = 28'b0000011000100110000011000000;
expected_data = 28'b0010110000000000000000000000;
@(next_data);

send_data = 28'b0001100101011000100100000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b1110001100101010100101000000;
expected_data = 28'b0011001000000000000000000000;
@(next_data);

send_data = 28'b0011011100110010000110000000;
expected_data = 28'b1001001001000000000000000000;
@(next_data);

send_data = 28'b1010001101101101000111000000;
expected_data = 28'b0011011100000000000000000000;
@(next_data);

send_data = 28'b1010010000111000001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0101000001111110101001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1011001001001010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010110001111111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1001011000111011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100011000001101001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110000010110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110101101001001001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011101011101100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011111000101010000001000000;
expected_data = 28'b1100001001000000000000000000;
@(next_data);

send_data = 28'b1111001001100111100010000000;
expected_data = 28'b0110101000000000000000000000;
@(next_data);

send_data = 28'b1110011000100011000011000000;
expected_data = 28'b1100001001000000000000000000;
@(next_data);

send_data = 28'b0111010100101000000100000000;
expected_data = 28'b0111001100000000000000000000;
@(next_data);

send_data = 28'b0001010001001101100101000000;
expected_data = 28'b1110101001000000000000000000;
@(next_data);

send_data = 28'b0111101100001101100110000000;
expected_data = 28'b0001111000000000000000000000;
@(next_data);

send_data = 28'b1100101000011100100111000000;
expected_data = 28'b0111101100000000000000000000;
@(next_data);

send_data = 28'b1010100101001011001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1010110001010100001001000000;
expected_data = 28'b0000100000100000000000000000;
@(next_data);

send_data = 28'b1000011000100101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0100001000110110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000011000100110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111010100110101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001010101010101001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010100100010000001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011010000111111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100101000100111000001000000;
expected_data = 28'b1011001001000000000000000000;
@(next_data);

send_data = 28'b1100011100000010100010000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0001111000000000000011000000;
expected_data = 28'b0011110100000000000000000000;
@(next_data);

send_data = 28'b0010011100101000000100000000;
expected_data = 28'b0000111100000000000000000000;
@(next_data);

send_data = 28'b0011101000101110000101000000;
expected_data = 28'b0100111000000000000000000000;
@(next_data);

send_data = 28'b0001001101101101000110000000;
expected_data = 28'b0010011100000000000000000000;
@(next_data);

send_data = 28'b1111010000100011100111000000;
expected_data = 28'b0001001100000000000000000000;
@(next_data);

send_data = 28'b1001000001011001001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1010001100100100001001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1110001100111110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1000100101010110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1010001101110110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011111000101100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000100001001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011100100001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100001100001000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111101100010010000001000000;
expected_data = 28'b0101001100000000000000000000;
@(next_data);

send_data = 28'b0011111000111110100010000000;
expected_data = 28'b0101111100000000000000000000;
@(next_data);

send_data = 28'b0010010100010100000011000000;
expected_data = 28'b1011110001000000000000000000;
@(next_data);

send_data = 28'b1001000000100001100100000000;
expected_data = 28'b0001001000000000000000000000;
@(next_data);

send_data = 28'b1100011000100011000101000000;
expected_data = 28'b0010000000100000000000000000;
@(next_data);

send_data = 28'b1001000100000011100110000000;
expected_data = 28'b1010010101000000000000000000;
@(next_data);

send_data = 28'b1011111100001111000111000000;
expected_data = 28'b1110111101000000000000000000;
@(next_data);

send_data = 28'b1101000001111001101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0010111001101101001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1101000100001000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1000010100000011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1011011101110001101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110000101110100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101110101000101101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111110100011010001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001011100001100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010001010110100001000000;
expected_data = 28'b0011000000000000000000000000;
@(next_data);

send_data = 28'b1000110000101011000010000000;
expected_data = 28'b1011100101000000000000000000;
@(next_data);

send_data = 28'b1000110001010010000011000000;
expected_data = 28'b0010010100000000000000000000;
@(next_data);

send_data = 28'b1110100001010111100100000000;
expected_data = 28'b0100011000000000000000000000;
@(next_data);

send_data = 28'b1100011001011111000101000000;
expected_data = 28'b1101000001000000000000000000;
@(next_data);

send_data = 28'b1110001001000000000110000000;
expected_data = 28'b1010010101000000000000000000;
@(next_data);

send_data = 28'b1110001000001010000111000000;
expected_data = 28'b1001111001000000000000000000;
@(next_data);

send_data = 28'b1011011000111111001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101111000000111101001000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1011001000110010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101000101111110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0110011001011010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011010101101111101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001001001010110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000000000110001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110100000011110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111010100111101000001000000;
expected_data = 28'b1010010101000000000000000000;
@(next_data);

send_data = 28'b0011110100010101000010000000;
expected_data = 28'b1000111101000000000000000000;
@(next_data);

send_data = 28'b1111110001001001000011000000;
expected_data = 28'b1110100001000000000000000000;
@(next_data);

send_data = 28'b0011111000001010000100000000;
expected_data = 28'b0111111000000000000000000000;
@(next_data);

send_data = 28'b1101101101110000100101000000;
expected_data = 28'b0111110000000000000000000000;
@(next_data);

send_data = 28'b0100011101001110100110000000;
expected_data = 28'b1011011001000000000000000000;
@(next_data);

send_data = 28'b0010101101011011000111000000;
expected_data = 28'b0100011100000000000000000000;
@(next_data);

send_data = 28'b0110100000111000101000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1101110000101010001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0011110100100110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010001100100101001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1010110101101110001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101001011010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111001000101001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100100111100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100101000001010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001000101101000000001000000;
expected_data = 28'b1101111101000000000000000000;
@(next_data);

send_data = 28'b0011011100000101000010000000;
expected_data = 28'b0100000100000000000000000000;
@(next_data);

send_data = 28'b0011001100100101000011000000;
expected_data = 28'b1100001001000000000000000000;
@(next_data);

send_data = 28'b0111101001110101000100000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b0100000101000011000101000000;
expected_data = 28'b1111010001000000000000000000;
@(next_data);

send_data = 28'b0101101100010111000110000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b1000000001100011000111000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b1110001101110001001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110101001100110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1000010000001011101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0100011101110000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0101111001100110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100011001001101101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100011101010111001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111100100101001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010010100011001100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011101011000100001000000;
expected_data = 28'b1101100001000000000000000000;
@(next_data);

send_data = 28'b1011010100111111100010000000;
expected_data = 28'b0100011000000000000000000000;
@(next_data);

send_data = 28'b0000101100101101000011000000;
expected_data = 28'b0011010100000000000000000000;
@(next_data);

send_data = 28'b0101110001010001000100000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b1100101100011100000101000000;
expected_data = 28'b1011100001000000000000000000;
@(next_data);

send_data = 28'b0001000100111100000110000000;
expected_data = 28'b1010111001000000000000000000;
@(next_data);

send_data = 28'b1101111100100001100111000000;
expected_data = 28'b0001000100000000000000000000;
@(next_data);

send_data = 28'b1111111001110000001000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b0110000100101001101001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1110111101000011101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0001111101110101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0010011001111010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100100111110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010110000001110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110110100000111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101100010000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100101101101001000001000000;
expected_data = 28'b0101110000000000000000000000;
@(next_data);

send_data = 28'b0100110101000101000010000000;
expected_data = 28'b0001100100000000000000000000;
@(next_data);

send_data = 28'b0111001101000100000011000000;
expected_data = 28'b0011100000000000000000000000;
@(next_data);

send_data = 28'b0111101101010001100100000000;
expected_data = 28'b0011100100000000000000000000;
@(next_data);

send_data = 28'b1110010000011111100101000000;
expected_data = 28'b1111011001000000000000000000;
@(next_data);

send_data = 28'b1011001100011101000110000000;
expected_data = 28'b1001011001000000000000000000;
@(next_data);

send_data = 28'b0101111100110000100111000000;
expected_data = 28'b1100110101000000000000000000;
@(next_data);

send_data = 28'b0110011000110111101000000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011000100111101101001000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0011111101101101001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1010101001100101101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1000100001011011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000101001111100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100010000101000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101010001111100101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010011000110000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100101001010010100001000000;
expected_data = 28'b0000011100010000000000000000;
@(next_data);

send_data = 28'b1110101101010001100010000000;
expected_data = 28'b1110111101000000000000000000;
@(next_data);

send_data = 28'b0111010101101001000011000000;
expected_data = 28'b1011011101000000000000000000;
@(next_data);

send_data = 28'b0100011100100110100100000000;
expected_data = 28'b0011101000000000000000000000;
@(next_data);

send_data = 28'b1001000001001011100101000000;
expected_data = 28'b1000111001000000000000000000;
@(next_data);

send_data = 28'b1110010101010110000110000000;
expected_data = 28'b1101100001000000000000000000;
@(next_data);

send_data = 28'b0010110101000101100111000000;
expected_data = 28'b1001101101000000000000000000;
@(next_data);

send_data = 28'b1010000001000111001000000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110010001001000101001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1000110001100010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1111101000001110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1101111100111000001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011100000110100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101111000011110101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110101001001110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101011100110110100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100101000100111100001000000;
expected_data = 28'b0100010000010000000000000000;
@(next_data);

send_data = 28'b1101010001011101100010000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0010111100110111100011000000;
expected_data = 28'b1001000001000000000000000000;
@(next_data);

send_data = 28'b0000011101111100100100000000;
expected_data = 28'b0001011100000000000000000000;
@(next_data);

send_data = 28'b0110101001111011000101000000;
expected_data = 28'b0000111000000000000000000000;
@(next_data);

send_data = 28'b1010000000111110100110000000;
expected_data = 28'b0101111100000000000000000000;
@(next_data);

send_data = 28'b1001000000110011100111000000;
expected_data = 28'b1110000001000000000000000000;
@(next_data);

send_data = 28'b0000101100011001101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001110001001100001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0100100000111010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0011110001011001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0110000100111001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001101001110000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001111100100110001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000101011100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001100001011011000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011011101011000100001000000;
expected_data = 28'b0100111000010000000000000000;
@(next_data);

send_data = 28'b1010010000011110000010000000;
expected_data = 28'b1000011001000000000000000000;
@(next_data);

send_data = 28'b1101101101100111000011000000;
expected_data = 28'b0110011100000000000000000000;
@(next_data);

send_data = 28'b1101110001111010100100000000;
expected_data = 28'b0110110100000000000000000000;
@(next_data);

send_data = 28'b1010010101100100100101000000;
expected_data = 28'b1011100001000000000000000000;
@(next_data);

send_data = 28'b0011011101101001100110000000;
expected_data = 28'b1111011101000000000000000000;
@(next_data);

send_data = 28'b1110011001101000000111000000;
expected_data = 28'b0011011100000000000000000000;
@(next_data);

send_data = 28'b1101101100100110001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000100100101101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011101001001000001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011010101001010001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0001011100000101101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011000000010100001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100000110000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000010000100010001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110001010011100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001100000110001000001000000;
expected_data = 28'b0011001100010000000000000000;
@(next_data);

send_data = 28'b0101000100000011100010000000;
expected_data = 28'b0111101000000000000000000000;
@(next_data);

send_data = 28'b1100011101001010100011000000;
expected_data = 28'b1010100101000000000000000000;
@(next_data);

send_data = 28'b1011110101000101100100000000;
expected_data = 28'b0110001100000000000000000000;
@(next_data);

send_data = 28'b0000101100011010100101000000;
expected_data = 28'b0111101000000000000000000000;
@(next_data);

send_data = 28'b0101011000100111000110000000;
expected_data = 28'b0000111000000000000000000000;
@(next_data);

send_data = 28'b1010010101101110000111000000;
expected_data = 28'b0101011000000000000000000000;
@(next_data);

send_data = 28'b0010000001011111001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1001010100001111001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1000010000011000101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1100000000000011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110011000111110101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001000001100000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110111001101011101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111001100111001001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010101101010001000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100101011000100001000000;
expected_data = 28'b1100110101000000000000000000;
@(next_data);

send_data = 28'b0010011100111010000010000000;
expected_data = 28'b0011100000000000000000000000;
@(next_data);

send_data = 28'b0101111001010001000011000000;
expected_data = 28'b1010110001000000000000000000;
@(next_data);

send_data = 28'b0111101001111100100100000000;
expected_data = 28'b0010111100000000000000000000;
@(next_data);

send_data = 28'b0000000100001100000101000000;
expected_data = 28'b1111010001000000000000000000;
@(next_data);

send_data = 28'b1111111100000010000110000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b0101101101101011000111000000;
expected_data = 28'b1000000101000000000000000000;
@(next_data);

send_data = 28'b1011111000110100001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0001000000011110001001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1001111101110111001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101001001000001101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1000101000000010101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110101001110010001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000001000000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110101001010101001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100011100000000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011111101010011100001000000;
expected_data = 28'b1100100001000000000000000000;
@(next_data);

send_data = 28'b1100101000101010000010000000;
expected_data = 28'b0001100000000000000000000000;
@(next_data);

send_data = 28'b0001111000000101100011000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b1011101000111100000100000000;
expected_data = 28'b0000111100000000000000000000;
@(next_data);

send_data = 28'b1000000100000100000101000000;
expected_data = 28'b0111010000000000000000000000;
@(next_data);

send_data = 28'b1000110001000010000110000000;
expected_data = 28'b1100000101000000000000000000;
@(next_data);

send_data = 28'b1010111100100001100111000000;
expected_data = 28'b1111010001000000000000000000;
@(next_data);

send_data = 28'b0111001100010000001000000000;
expected_data = 28'b0000000100100000000000000000;
@(next_data);

send_data = 28'b0000010101000100001001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b0101101001101001101010000000;
expected_data = 28'b0001111100000000000000000000;
@(next_data);

send_data = 28'b0111011001011110101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1001011101101011101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000011001000010001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100010101010100101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001101001000110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000101000001010100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000100000000000100001000000;
expected_data = 28'b1001111101000000000000000000;
@(next_data);

send_data = 28'b0011100001111000000010000000;
expected_data = 28'b1000100101000000000000000000;
@(next_data);

send_data = 28'b1010000000010000000011000000;
expected_data = 28'b0011011100000000000000000000;
@(next_data);

send_data = 28'b1111110100011100000100000000;
expected_data = 28'b0101000000000000000000000000;
@(next_data);

send_data = 28'b0001111100101001000101000000;
expected_data = 28'b1111101001000000000000000000;
@(next_data);

send_data = 28'b1011000101101010100110000000;
expected_data = 28'b0001000000100000000000000000;
@(next_data);

send_data = 28'b0101111001110000000111000000;
expected_data = 28'b1100111101000000000000000000;
@(next_data);

send_data = 28'b1101010001011001101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110001001111101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110000000110011101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0101001001001111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0111011100001111101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100000100100100101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1001110000001001101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100111101111000001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111011000010100100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0100100100011100000001000000;
expected_data = 28'b1001111101000000000000000000;
@(next_data);

send_data = 28'b1100010000000101000010000000;
expected_data = 28'b0111000100000000000000000000;
@(next_data);

send_data = 28'b1001010000110011000011000000;
expected_data = 28'b0011000100000000000000000000;
@(next_data);

send_data = 28'b1001101100110000100100000000;
expected_data = 28'b0100101000000000000000000000;
@(next_data);

send_data = 28'b0000011001111101100101000000;
expected_data = 28'b0011011000000000000000000000;
@(next_data);

send_data = 28'b0111100000111011100110000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0100000001010000100111000000;
expected_data = 28'b0111100000000000000000000000;
@(next_data);

send_data = 28'b0101000101110100001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101011001101001001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1010111101010010101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0010000100100100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0110111000000000101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010001001011001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011101101111101001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110100101110100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110010000111111000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111111100111110000001000000;
expected_data = 28'b1110001001000000000000000000;
@(next_data);

send_data = 28'b0001110101101100100010000000;
expected_data = 28'b1000001101000000000000000000;
@(next_data);

send_data = 28'b1100001101001110000011000000;
expected_data = 28'b0011101100000000000000000000;
@(next_data);

send_data = 28'b1100001100001001000100000000;
expected_data = 28'b0110000100000000000000000000;
@(next_data);

send_data = 28'b1111100101100000100101000000;
expected_data = 28'b1000011001000000000000000000;
@(next_data);

send_data = 28'b0100001100101111100110000000;
expected_data = 28'b1000010101000000000000000000;
@(next_data);

send_data = 28'b0100001001011001000111000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b0010110100111110001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1010110000010111101001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1010001000000001001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1011011100001100001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1001101001001100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1000110101000001101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011000100001000001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110001101011110001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000011000100111100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011111101011001100001000000;
expected_data = 28'b0101010100000000000000000000;
@(next_data);

send_data = 28'b0100011000001000000010000000;
expected_data = 28'b1000110001000000000000000000;
@(next_data);

send_data = 28'b0000110001011100100011000000;
expected_data = 28'b1010100101000000000000000000;
@(next_data);

send_data = 28'b0111111000110010000100000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0101001100001100100101000000;
expected_data = 28'b1111110001000000000000000000;
@(next_data);

send_data = 28'b1100110101111111000110000000;
expected_data = 28'b0111101000000000000000000000;
@(next_data);

send_data = 28'b0110100100111100000111000000;
expected_data = 28'b1011001101000000000000000000;
@(next_data);

send_data = 28'b1000011100010010101000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0111000100111100001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1110100000110110001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0000000101001111001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1110110001111100001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101010101110000101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110010101000000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0101000001110101101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110011001100110000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0011011000111110100001000000;
expected_data = 28'b1011001001010000000000000000;
@(next_data);

send_data = 28'b1001110001101011100010000000;
expected_data = 28'b0100101100000000000000000000;
@(next_data);

send_data = 28'b0110011101110101100011000000;
expected_data = 28'b1011010001000000000000000000;
@(next_data);

send_data = 28'b1010101100110011000100000000;
expected_data = 28'b0011001100000000000000000000;
@(next_data);

send_data = 28'b0000011100011000100101000000;
expected_data = 28'b0101011000000000000000000000;
@(next_data);

send_data = 28'b0010101000011101000110000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1101011001000111100111000000;
expected_data = 28'b0010101000000000000000000000;
@(next_data);

send_data = 28'b0101010101001001001000000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b0001110000010100101001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b0000101100100100001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b0000001001010011001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0011000000010111101100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010100100011110001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001010101111000001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101101000010111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110010100010001000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101000011000100001000000;
expected_data = 28'b1000011101000000000000000000;
@(next_data);

send_data = 28'b1101001101100111100010000000;
expected_data = 28'b1001101101000000000000000000;
@(next_data);

send_data = 28'b1110011001001100000011000000;
expected_data = 28'b1110001101000000000000000000;
@(next_data);

send_data = 28'b0000000100010001000100000000;
expected_data = 28'b0111001100000000000000000000;
@(next_data);

send_data = 28'b1010000101110111000101000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1100001100111001000110000000;
expected_data = 28'b1111000101000000000000000000;
@(next_data);

send_data = 28'b1011110101100110000111000000;
expected_data = 28'b1011110101000000000000000000;
@(next_data);

send_data = 28'b0110010000110100001000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b1011111100111010101001000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1110101000111001001010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1101100000011000001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0000110000011111001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110000101101001001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101100000111011001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1100001000111100001111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1011110100111000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1111011101110000000001000000;
expected_data = 28'b0010110100010000000000000000;
@(next_data);

send_data = 28'b1111101000001000000010000000;
expected_data = 28'b0001011100000000000000000000;
@(next_data);

send_data = 28'b1010111100101111100011000000;
expected_data = 28'b0001010100000000000000000000;
@(next_data);

send_data = 28'b0001000001001010100100000000;
expected_data = 28'b0101011100000000000000000000;
@(next_data);

send_data = 28'b0100010001110111000101000000;
expected_data = 28'b0010000000100000000000000000;
@(next_data);

send_data = 28'b0101101100111110000110000000;
expected_data = 28'b0110011000000000000000000000;
@(next_data);

send_data = 28'b0110110100011101100111000000;
expected_data = 28'b0101101100000000000000000000;
@(next_data);

send_data = 28'b0101101000100010101000000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0000010000100100001001000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1100000000011111101010000000;
expected_data = 28'b0000111100000000000000000000;
@(next_data);

send_data = 28'b1011010100111100101011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b1111100100010010001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110110101010000001101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001110001010100001110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1110001101110111101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0000000001101000100000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0001001100101000000001000000;
expected_data = 28'b1101000101000000000000000000;
@(next_data);

send_data = 28'b0111001100010110100010000000;
expected_data = 28'b0100001100000000000000000000;
@(next_data);

send_data = 28'b0000010000001011000011000000;
expected_data = 28'b1010000101000000000000000000;
@(next_data);

send_data = 28'b0100000001011100100100000000;
expected_data = 28'b0000001000100000000000000000;
@(next_data);

send_data = 28'b1010101101000010100101000000;
expected_data = 28'b1000000001100000000000000000;
@(next_data);

send_data = 28'b0000111001010100000110000000;
expected_data = 28'b1111111001000000000000000000;
@(next_data);

send_data = 28'b0100110000010000100111000000;
expected_data = 28'b0000111000000000000000000000;
@(next_data);

send_data = 28'b1011010001011111101000000000;
expected_data = 28'b0000010000100000000000000000;
@(next_data);

send_data = 28'b0010101100100010101001000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0001110000111110101010000000;
expected_data = 28'b1111111111010000000000000000;
@(next_data);

send_data = 28'b1110011101111001001011000000;
expected_data = 28'b0000000000010000000000000000;
@(next_data);

send_data = 28'b0100110001101001001100000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1101001100101010101101000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010101001001000101110000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0010111101111001101111000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);
